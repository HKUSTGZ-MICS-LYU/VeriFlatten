module fpu (
	clk,
	rmode,
	fpu_op,
	opa,
	opb,
	sender_valid,
	out,
	inf,
	snan,
	qnan,
	ine,
	overflow,
	underflow,
	zero,
	div_by_zero,
	input_ready,
	output_valid
);
	reg [31:0] ___sel_temp_0;
	reg [31:0] ___sel_temp_1;
	reg [31:0] ___sel_temp_2;
	reg [31:0] ___sel_temp_3;
	wire [8:0] ___sel_temp_4;
	wire [8:0] ___sel_temp_5;
	wire [8:0] ___sel_temp_6;
	wire [8:0] ___sel_temp_7;
	wire [31:0] ___sel_temp_8;
	wire [27:0] ___sel_temp_9;
	wire [27:0] ___sel_temp_10;
	wire [24:0] ___sel_temp_11;
	wire [24:0] ___sel_temp_12;
	wire [24:0] ___sel_temp_13;
	wire [24:0] ___sel_temp_14;
	wire [24:0] ___sel_temp_15;
	wire [24:0] ___sel_temp_16;
	wire [24:0] ___sel_temp_17;
	wire [24:0] ___sel_temp_18;
	wire [24:0] ___sel_temp_19;
	wire [24:0] ___sel_temp_20;
	wire [24:0] ___sel_temp_21;
	wire [24:0] ___sel_temp_22;
	wire [24:0] ___sel_temp_23;
	wire [24:0] ___sel_temp_24;
	wire [24:0] ___sel_temp_25;
	wire [24:0] ___sel_temp_26;
	wire [24:0] ___sel_temp_27;
	wire [24:0] ___sel_temp_28;
	wire [24:0] ___sel_temp_29;
	wire [24:0] ___sel_temp_30;
	wire [24:0] ___sel_temp_31;
	wire [24:0] ___sel_temp_32;
	wire [24:0] ___sel_temp_33;
	wire [24:0] ___sel_temp_34;
	wire [24:0] ___sel_temp_35;
	wire [24:0] ___sel_temp_36;
	wire [24:0] ___sel_temp_37;
	wire [24:0] ___sel_temp_38;
	wire [24:0] ___sel_temp_39;
	wire [24:0] ___sel_temp_40;
	wire [24:0] ___sel_temp_41;
	wire [24:0] ___sel_temp_42;
	wire [24:0] ___sel_temp_43;
	wire [24:0] ___sel_temp_44;
	wire [24:0] ___sel_temp_45;
	wire [24:0] ___sel_temp_46;
	wire [24:0] ___sel_temp_47;
	wire [24:0] ___sel_temp_48;
	wire [24:0] ___sel_temp_49;
	wire [24:0] ___sel_temp_50;
	wire [24:0] ___sel_temp_51;
	wire [24:0] ___sel_temp_52;
	wire [24:0] ___sel_temp_53;
	wire [24:0] ___sel_temp_54;
	wire [24:0] ___sel_temp_55;
	wire [24:0] ___sel_temp_56;
	wire [24:0] ___sel_temp_57;
	wire [24:0] ___sel_temp_58;
	wire [24:0] ___sel_temp_59;
	wire [24:0] ___sel_temp_60;
	wire [8:0] ___sel_temp_61;
	wire [8:0] ___sel_temp_62;
	wire [8:0] ___sel_temp_63;
	wire [8:0] ___sel_temp_64;
	wire [31:0] ___sel_temp_65;
	wire [31:0] ___sel_temp_66;
	wire [31:0] ___sel_temp_67;
	wire [47:0] ___sel_temp_68;
	wire [47:0] ___sel_temp_69;
	wire [8:0] ___sel_temp_70;
	wire [8:0] ___sel_temp_71;
	wire [31:0] ___sel_temp_72;
	wire [31:0] ___sel_temp_73;
	wire [31:0] ___sel_temp_74;
	wire [31:0] ___sel_temp_75;
	wire [23:0] ___sel_temp_76;
	wire [23:0] ___sel_temp_77;
	wire [23:0] ___sel_temp_78;
	wire [23:0] ___sel_temp_79;
	input wire clk;
	input wire [1:0] rmode;
	input wire [2:0] fpu_op;
	input wire [31:0] opa;
	input wire [31:0] opb;
	input wire sender_valid;
	output reg [31:0] out;
	output reg inf;
	output reg snan;
	output reg qnan;
	output reg ine;
	output reg overflow;
	output reg underflow;
	output reg zero;
	output reg div_by_zero;
	output reg input_ready;
	output reg output_valid;
	wire fpu___clk;
	wire [1:0] fpu___rmode;
	wire [2:0] fpu___fpu_op;
	wire [31:0] fpu___opa;
	wire [31:0] fpu___opb;
	wire fpu___sender_valid;
	reg [31:0] fpu___out;
	reg fpu___inf;
	reg fpu___snan;
	reg fpu___qnan;
	reg fpu___ine;
	reg fpu___overflow;
	reg fpu___underflow;
	reg fpu___zero;
	reg fpu___div_by_zero;
	reg fpu___input_ready;
	reg fpu___output_valid;
	parameter [30:0] fpu___INF = 31'h7f800000;
	parameter [30:0] fpu___QNAN = 31'h7fc00001;
	parameter [30:0] fpu___SNAN = 31'h7f800001;
	reg fpu___data_accept_r1;
	reg fpu___data_accept_r2;
	reg fpu___data_accept_r3;
	reg [31:0] fpu___opa_r;
	reg [31:0] fpu___opb_r;
	wire fpu___signa;
	wire fpu___signb;
	reg fpu___sign_fasu;
	reg [26:0] fpu___fracta;
	reg [26:0] fpu___fractb;
	reg [7:0] fpu___exp_fasu;
	reg [7:0] fpu___exp_r;
	wire [26:0] fpu___fract_out_d;
	wire fpu___co;
	reg [27:0] fpu___fract_out_q;
	wire [30:0] fpu___out_d;
	wire fpu___overflow_d;
	wire fpu___underflow_d;
	reg [1:0] fpu___rmode_r1;
	reg [1:0] fpu___rmode_r2;
	reg [1:0] fpu___rmode_r3;
	reg [2:0] fpu___fpu_op_r1;
	reg [2:0] fpu___fpu_op_r2;
	reg [2:0] fpu___fpu_op_r3;
	wire fpu___mul_inf;
	wire fpu___div_inf;
	wire fpu___mul_00;
	wire fpu___div_00;
	reg fpu___inf_d;
	reg fpu___ind_d;
	reg fpu___qnan_d;
	reg fpu___snan_d;
	reg fpu___opa_nan;
	reg fpu___opb_nan;
	reg fpu___opa_00;
	reg fpu___opb_00;
	reg fpu___opa_inf;
	reg fpu___opb_inf;
	reg fpu___opa_dn;
	reg fpu___opb_dn;
	reg fpu___nan_sign_d;
	reg fpu___result_zero_sign_d;
	reg fpu___sign_fasu_r;
	reg [7:0] fpu___exp_mul;
	reg fpu___sign_mul;
	reg fpu___sign_mul_r;
	wire [23:0] fpu___fracta_mul;
	wire [23:0] fpu___fractb_mul;
	reg fpu___inf_mul;
	reg fpu___inf_mul_r;
	reg [1:0] fpu___exp_ovf;
	reg [1:0] fpu___exp_ovf_r;
	reg fpu___sign_exe;
	reg fpu___sign_exe_r;
	reg [2:0] fpu___underflow_fmul_d;
	wire fpu_____Vcellinp__u1__add;
	reg [47:0] fpu___prod;
	wire [49:0] fpu___quo;
	wire [49:0] fpu___fdiv_opa;
	wire [49:0] fpu___remainder;
	wire fpu___remainder_00;
	reg [4:0] fpu___div_opa_ldz_d;
	reg [4:0] fpu___div_opa_ldz_r1;
	reg [4:0] fpu___div_opa_ldz_r2;
	wire [23:0] fpu_____Vcellout__u_divider__remainder;
	wire fpu___ine_d;
	reg [47:0] fpu___fract_denorm;
	wire [47:0] fpu___fract_div;
	wire fpu___sign_d;
	reg fpu___sign;
	reg [30:0] fpu___opa_r1;
	reg [47:0] fpu___fract_i2f;
	reg fpu___opas_r1;
	reg fpu___opas_r2;
	wire fpu___f2i_out_sign;
	wire fpu_____Vcellinp__u4__output_zero;
	reg fpu___fasu_op_r1;
	reg fpu___fasu_op_r2;
	wire [30:0] fpu___out_fixed;
	wire fpu___output_zero_fasu;
	wire fpu___output_zero_fdiv;
	wire fpu___output_zero_fmul;
	reg fpu___inf_mul2;
	wire fpu___overflow_fasu;
	wire fpu___overflow_fmul;
	wire fpu___overflow_fdiv;
	wire fpu___inf_fmul;
	wire fpu___sign_mul_final;
	wire fpu___out_d_00;
	wire fpu___sign_div_final;
	wire fpu___ine_mul;
	wire fpu___ine_mula;
	wire fpu___ine_div;
	wire fpu___ine_fasu;
	wire fpu___underflow_fasu;
	wire fpu___underflow_fmul;
	wire fpu___underflow_fdiv;
	wire fpu___underflow_fmul1;
	reg [2:0] fpu___underflow_fmul_r;
	reg fpu___opa_nan_r;
	reg fpu___fasu_op;
	wire fpu___co_d;
	wire fpu___u0___clk;
	wire [31:0] fpu___u0___opa;
	wire [31:0] fpu___u0___opb;
	reg fpu___u0___inf;
	reg fpu___u0___ind;
	reg fpu___u0___qnan;
	reg fpu___u0___snan;
	reg fpu___u0___opa_nan;
	reg fpu___u0___opb_nan;
	reg fpu___u0___opa_00;
	reg fpu___u0___opb_00;
	reg fpu___u0___opa_inf;
	reg fpu___u0___opb_inf;
	reg fpu___u0___opa_dn;
	reg fpu___u0___opb_dn;
	wire [7:0] fpu___u0___expa;
	wire [7:0] fpu___u0___expb;
	wire [22:0] fpu___u0___fracta;
	wire [22:0] fpu___u0___fractb;
	reg fpu___u0___expa_ff;
	reg fpu___u0___infa_f_r;
	reg fpu___u0___qnan_r_a;
	reg fpu___u0___snan_r_a;
	reg fpu___u0___expb_ff;
	reg fpu___u0___infb_f_r;
	reg fpu___u0___qnan_r_b;
	reg fpu___u0___snan_r_b;
	reg fpu___u0___expa_00;
	reg fpu___u0___expb_00;
	reg fpu___u0___fracta_00;
	reg fpu___u0___fractb_00;
	wire fpu___u1___clk;
	wire [1:0] fpu___u1___rmode;
	wire fpu___u1___add;
	wire [31:0] fpu___u1___opa;
	wire [31:0] fpu___u1___opb;
	wire fpu___u1___opa_nan;
	wire fpu___u1___opb_nan;
	reg [26:0] fpu___u1___fracta_out;
	reg [26:0] fpu___u1___fractb_out;
	reg [7:0] fpu___u1___exp_dn_out;
	reg fpu___u1___sign;
	reg fpu___u1___nan_sign;
	reg fpu___u1___result_zero_sign;
	reg fpu___u1___fasu_op;
	wire fpu___u1___signa;
	wire fpu___u1___signb;
	wire [7:0] fpu___u1___expa;
	wire [7:0] fpu___u1___expb;
	wire [22:0] fpu___u1___fracta;
	wire [22:0] fpu___u1___fractb;
	wire fpu___u1___expa_lt_expb;
	wire fpu___u1___fractb_lt_fracta;
	wire [7:0] fpu___u1___exp_small;
	wire [7:0] fpu___u1___exp_large;
	wire [7:0] fpu___u1___exp_diff;
	wire [22:0] fpu___u1___adj_op;
	wire [26:0] fpu___u1___adj_op_tmp;
	wire [26:0] fpu___u1___adj_op_out;
	wire [26:0] fpu___u1___fracta_n;
	wire [26:0] fpu___u1___fractb_n;
	wire [26:0] fpu___u1___fracta_s;
	wire [26:0] fpu___u1___fractb_s;
	reg fpu___u1___sign_d;
	reg fpu___u1___add_d;
	wire fpu___u1___expa_dn;
	wire fpu___u1___expb_dn;
	reg fpu___u1___sticky;
	reg fpu___u1___add_r;
	reg fpu___u1___signa_r;
	reg fpu___u1___signb_r;
	wire [4:0] fpu___u1___exp_diff_sft;
	wire fpu___u1___exp_lt_27;
	wire fpu___u1___op_dn;
	wire [26:0] fpu___u1___adj_op_out_sft;
	reg fpu___u1___fracta_lt_fractb;
	reg fpu___u1___fracta_eq_fractb;
	wire fpu___u1___nan_sign1;
	wire [7:0] fpu___u1___exp_diff1;
	wire [7:0] fpu___u1___exp_diff1a;
	wire [7:0] fpu___u1___exp_diff2;
	wire fpu___u2___clk;
	wire [2:0] fpu___u2___fpu_op;
	wire [31:0] fpu___u2___opa;
	wire [31:0] fpu___u2___opb;
	wire [23:0] fpu___u2___fracta;
	wire [23:0] fpu___u2___fractb;
	reg [7:0] fpu___u2___exp_out;
	reg fpu___u2___sign;
	reg fpu___u2___sign_exe;
	reg fpu___u2___inf;
	reg [1:0] fpu___u2___exp_ovf;
	reg [2:0] fpu___u2___underflow;
	wire fpu___u2___signa;
	wire fpu___u2___signb;
	reg fpu___u2___sign_d;
	wire [1:0] fpu___u2___exp_ovf_d;
	wire [7:0] fpu___u2___expa;
	wire [7:0] fpu___u2___expb;
	wire [7:0] fpu___u2___exp_tmp1;
	wire [7:0] fpu___u2___exp_tmp2;
	wire fpu___u2___co1;
	wire fpu___u2___co2;
	wire fpu___u2___expa_dn;
	wire fpu___u2___expb_dn;
	wire [7:0] fpu___u2___exp_out_a;
	wire fpu___u2___opa_00;
	wire fpu___u2___opb_00;
	wire fpu___u2___fracta_00;
	wire fpu___u2___fractb_00;
	wire [7:0] fpu___u2___exp_tmp3;
	wire [7:0] fpu___u2___exp_tmp4;
	wire [7:0] fpu___u2___exp_tmp5;
	wire [2:0] fpu___u2___underflow_d;
	wire fpu___u2___op_div;
	wire [7:0] fpu___u2___exp_out_mul;
	wire [7:0] fpu___u2___exp_out_div;
	wire fpu___u3___add;
	wire [26:0] fpu___u3___opa;
	wire [26:0] fpu___u3___opb;
	wire [26:0] fpu___u3___sum;
	wire fpu___u3___co;
	wire fpu___u5___clk;
	wire [23:0] fpu___u5___opa;
	wire [23:0] fpu___u5___opb;
	reg [47:0] fpu___u5___prod;
	reg [47:0] fpu___u5___prod1;
	parameter [31:0] fpu___u_divider___N = 32'sh00000032;
	parameter [31:0] fpu___u_divider___M = 32'sh00000018;
	parameter [31:0] fpu___u_divider___N_ACT = 32'h00000049;
	parameter [31:0] fpu___u_divider___N_ACT_M = 32'h00000031;
	parameter [31:0] fpu___u_divider___PART1 = 32'h00000010;
	parameter [31:0] fpu___u_divider___PART2 = 32'h00000010;
	parameter [31:0] fpu___u_divider___PART3 = 32'h00000011;
	wire fpu___u_divider___clk;
	wire [49:0] fpu___u_divider___dividend;
	wire [23:0] fpu___u_divider___divisor;
	wire [49:0] fpu___u_divider___merchant;
	wire [23:0] fpu___u_divider___remainder;
	wire [48:0] fpu___u_divider___dividend_t1 [16:0];
	wire [23:0] fpu___u_divider___divisor_t1 [16:0];
	wire [49:0] fpu___u_divider___merchant_t1 [16:0];
	wire [23:0] fpu___u_divider___remainder_t1 [16:0];
	wire [48:0] fpu___u_divider___dividend_t2 [16:0];
	wire [23:0] fpu___u_divider___divisor_t2 [16:0];
	wire [49:0] fpu___u_divider___merchant_t2 [16:0];
	wire [23:0] fpu___u_divider___remainder_t2 [16:0];
	wire [48:0] fpu___u_divider___dividend_t3 [17:0];
	wire [23:0] fpu___u_divider___divisor_t3 [17:0];
	wire [49:0] fpu___u_divider___merchant_t3 [17:0];
	wire [23:0] fpu___u_divider___remainder_t3 [17:0];
	wire [23:0] fpu___u_divider_____Vcellout__u_divider_step0__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__u_divider_step0__merchant;
	wire [23:0] fpu___u_divider_____Vcellout__u_divider_step0__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellout__u_divider_step0__dividend_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__u_divider_step0__dividend_ci;
	wire [24:0] fpu___u_divider_____Vcellinp__u_divider_step0__dividend;
	reg [48:0] fpu___u_divider___dividend_t2_r;
	reg [23:0] fpu___u_divider___divisor_t2_r;
	reg [49:0] fpu___u_divider___merchant_t2_r;
	reg [23:0] fpu___u_divider___remainder_t2_r;
	reg [48:0] fpu___u_divider___dividend_t3_r;
	reg [23:0] fpu___u_divider___divisor_t3_r;
	reg [49:0] fpu___u_divider___merchant_t3_r;
	reg [23:0] fpu___u_divider___remainder_t3_r;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__remainder;
	wire [49:0] fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__merchant;
	wire [48:0] fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__dividend_kp;
	wire [23:0] fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__divisor_kp;
	wire [48:0] fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend_ci;
	wire [49:0] fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__merchant_ci;
	wire [23:0] fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__divisor;
	wire [24:0] fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend;
	parameter [31:0] fpu___u_divider___u_divider_step0___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___u_divider_step0___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___u_divider_step0___dividend;
	wire [23:0] fpu___u_divider___u_divider_step0___divisor;
	reg [49:0] fpu___u_divider___u_divider_step0___merchant_ci;
	initial fpu___u_divider___u_divider_step0___merchant_ci = 50'h0000000000000;
	wire [48:0] fpu___u_divider___u_divider_step0___dividend_ci;
	wire [48:0] fpu___u_divider___u_divider_step0___dividend_kp;
	wire [23:0] fpu___u_divider___u_divider_step0___divisor_kp;
	wire [49:0] fpu___u_divider___u_divider_step0___merchant;
	wire [23:0] fpu___u_divider___u_divider_step0___remainder;
	wire fpu___u_divider___u_divider_step0___geq;
	parameter [31:0] fpu___u_divider___gen_part11___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part11___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part11___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part11___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part11___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part11___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part11___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part11___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part11___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part11___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part11___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part12___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part12___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part12___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part12___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part12___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part12___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part12___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part12___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part12___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part12___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part12___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part13___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part13___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part13___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part13___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part13___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part13___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part13___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part13___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part13___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part13___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part13___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part14___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part14___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part14___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part14___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part14___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part14___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part14___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part14___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part14___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part14___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part14___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part15___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part15___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part15___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part15___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part15___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part15___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part15___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part15___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part15___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part15___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part15___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part16___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part16___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part16___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part16___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part16___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part16___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part16___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part16___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part16___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part16___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part16___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part17___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part17___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part17___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part17___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part17___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part17___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part17___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part17___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part17___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part17___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part17___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part18___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part18___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part18___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part18___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part18___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part18___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part18___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part18___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part18___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part18___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part18___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part19___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part19___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part19___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part19___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part19___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part19___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part19___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part19___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part19___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part19___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part19___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part110___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part110___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part110___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part110___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part110___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part110___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part110___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part110___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part110___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part110___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part110___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part111___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part111___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part111___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part111___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part111___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part111___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part111___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part111___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part111___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part111___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part111___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part112___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part112___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part112___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part112___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part112___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part112___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part112___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part112___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part112___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part112___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part112___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part113___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part113___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part113___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part113___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part113___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part113___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part113___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part113___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part113___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part113___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part113___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part114___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part114___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part114___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part114___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part114___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part114___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part114___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part114___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part114___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part114___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part114___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part115___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part115___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part115___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part115___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part115___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part115___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part115___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part115___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part115___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part115___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part115___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part116___u_divider_step1___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part116___u_divider_step1___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part116___u_divider_step1___dividend;
	wire [23:0] fpu___u_divider___gen_part116___u_divider_step1___divisor;
	wire [49:0] fpu___u_divider___gen_part116___u_divider_step1___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part116___u_divider_step1___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part116___u_divider_step1___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part116___u_divider_step1___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part116___u_divider_step1___merchant;
	wire [23:0] fpu___u_divider___gen_part116___u_divider_step1___remainder;
	wire fpu___u_divider___gen_part116___u_divider_step1___geq;
	parameter [31:0] fpu___u_divider___gen_part21___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part21___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part21___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part21___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part21___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part21___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part21___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part21___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part21___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part21___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part21___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part22___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part22___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part22___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part22___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part22___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part22___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part22___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part22___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part22___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part22___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part22___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part23___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part23___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part23___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part23___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part23___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part23___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part23___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part23___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part23___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part23___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part23___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part24___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part24___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part24___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part24___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part24___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part24___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part24___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part24___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part24___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part24___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part24___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part25___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part25___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part25___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part25___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part25___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part25___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part25___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part25___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part25___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part25___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part25___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part26___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part26___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part26___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part26___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part26___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part26___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part26___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part26___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part26___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part26___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part26___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part27___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part27___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part27___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part27___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part27___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part27___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part27___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part27___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part27___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part27___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part27___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part28___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part28___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part28___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part28___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part28___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part28___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part28___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part28___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part28___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part28___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part28___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part29___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part29___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part29___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part29___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part29___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part29___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part29___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part29___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part29___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part29___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part29___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part210___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part210___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part210___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part210___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part210___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part210___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part210___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part210___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part210___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part210___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part210___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part211___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part211___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part211___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part211___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part211___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part211___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part211___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part211___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part211___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part211___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part211___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part212___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part212___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part212___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part212___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part212___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part212___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part212___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part212___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part212___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part212___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part212___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part213___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part213___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part213___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part213___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part213___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part213___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part213___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part213___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part213___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part213___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part213___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part214___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part214___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part214___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part214___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part214___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part214___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part214___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part214___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part214___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part214___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part214___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part215___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part215___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part215___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part215___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part215___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part215___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part215___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part215___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part215___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part215___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part215___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part216___u_divider_step2___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part216___u_divider_step2___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part216___u_divider_step2___dividend;
	wire [23:0] fpu___u_divider___gen_part216___u_divider_step2___divisor;
	wire [49:0] fpu___u_divider___gen_part216___u_divider_step2___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part216___u_divider_step2___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part216___u_divider_step2___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part216___u_divider_step2___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part216___u_divider_step2___merchant;
	wire [23:0] fpu___u_divider___gen_part216___u_divider_step2___remainder;
	wire fpu___u_divider___gen_part216___u_divider_step2___geq;
	parameter [31:0] fpu___u_divider___gen_part31___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part31___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part31___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part31___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part31___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part31___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part31___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part31___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part31___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part31___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part31___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part32___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part32___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part32___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part32___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part32___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part32___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part32___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part32___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part32___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part32___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part32___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part33___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part33___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part33___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part33___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part33___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part33___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part33___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part33___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part33___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part33___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part33___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part34___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part34___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part34___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part34___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part34___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part34___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part34___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part34___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part34___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part34___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part34___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part35___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part35___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part35___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part35___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part35___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part35___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part35___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part35___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part35___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part35___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part35___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part36___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part36___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part36___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part36___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part36___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part36___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part36___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part36___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part36___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part36___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part36___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part37___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part37___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part37___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part37___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part37___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part37___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part37___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part37___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part37___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part37___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part37___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part38___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part38___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part38___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part38___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part38___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part38___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part38___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part38___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part38___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part38___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part38___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part39___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part39___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part39___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part39___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part39___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part39___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part39___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part39___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part39___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part39___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part39___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part310___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part310___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part310___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part310___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part310___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part310___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part310___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part310___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part310___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part310___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part310___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part311___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part311___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part311___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part311___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part311___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part311___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part311___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part311___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part311___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part311___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part311___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part312___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part312___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part312___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part312___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part312___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part312___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part312___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part312___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part312___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part312___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part312___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part313___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part313___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part313___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part313___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part313___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part313___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part313___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part313___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part313___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part313___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part313___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part314___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part314___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part314___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part314___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part314___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part314___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part314___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part314___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part314___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part314___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part314___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part315___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part315___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part315___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part315___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part315___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part315___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part315___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part315___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part315___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part315___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part315___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part316___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part316___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part316___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part316___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part316___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part316___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part316___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part316___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part316___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part316___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part316___u_divider_step3___geq;
	parameter [31:0] fpu___u_divider___gen_part317___u_divider_step3___N = 32'h00000049;
	parameter [31:0] fpu___u_divider___gen_part317___u_divider_step3___M = 32'sh00000018;
	wire [24:0] fpu___u_divider___gen_part317___u_divider_step3___dividend;
	wire [23:0] fpu___u_divider___gen_part317___u_divider_step3___divisor;
	wire [49:0] fpu___u_divider___gen_part317___u_divider_step3___merchant_ci;
	wire [48:0] fpu___u_divider___gen_part317___u_divider_step3___dividend_ci;
	wire [48:0] fpu___u_divider___gen_part317___u_divider_step3___dividend_kp;
	wire [23:0] fpu___u_divider___gen_part317___u_divider_step3___divisor_kp;
	wire [49:0] fpu___u_divider___gen_part317___u_divider_step3___merchant;
	wire [23:0] fpu___u_divider___gen_part317___u_divider_step3___remainder;
	wire fpu___u_divider___gen_part317___u_divider_step3___geq;
	wire fpu___u4___clk;
	wire [2:0] fpu___u4___fpu_op;
	wire fpu___u4___opas;
	wire fpu___u4___sign;
	wire [1:0] fpu___u4___rmode;
	wire [47:0] fpu___u4___fract_in;
	wire [7:0] fpu___u4___exp_in;
	wire [1:0] fpu___u4___exp_ovf;
	wire fpu___u4___opa_dn;
	wire fpu___u4___opb_dn;
	wire fpu___u4___rem_00;
	wire [4:0] fpu___u4___div_opa_ldz;
	wire fpu___u4___output_zero;
	wire [30:0] fpu___u4___out;
	wire fpu___u4___ine;
	wire fpu___u4___overflow;
	wire fpu___u4___underflow;
	wire fpu___u4___f2i_out_sign;
	wire [22:0] fpu___u4___fract_out;
	wire [7:0] fpu___u4___exp_out;
	wire fpu___u4___exp_out1_co;
	wire [22:0] fpu___u4___fract_out_final;
	reg [22:0] fpu___u4___fract_out_rnd;
	wire [8:0] fpu___u4___exp_next_mi;
	wire fpu___u4___dn;
	wire fpu___u4___exp_rnd_adj;
	wire [7:0] fpu___u4___exp_out_final;
	reg [7:0] fpu___u4___exp_out_rnd;
	wire fpu___u4___op_dn;
	wire fpu___u4___op_mul;
	wire fpu___u4___op_div;
	wire fpu___u4___op_i2f;
	wire fpu___u4___op_f2i;
	reg [5:0] fpu___u4___fi_ldz;
	wire fpu___u4___g;
	wire fpu___u4___r;
	wire fpu___u4___s;
	wire fpu___u4___round;
	wire fpu___u4___round2;
	wire fpu___u4___round2a;
	wire fpu___u4___round2_fasu;
	wire fpu___u4___round2_fmul;
	wire [7:0] fpu___u4___exp_out_rnd0;
	wire [7:0] fpu___u4___exp_out_rnd1;
	wire [7:0] fpu___u4___exp_out_rnd2;
	wire [7:0] fpu___u4___exp_out_rnd2a;
	wire [22:0] fpu___u4___fract_out_rnd0;
	wire [22:0] fpu___u4___fract_out_rnd1;
	wire [22:0] fpu___u4___fract_out_rnd2;
	wire [22:0] fpu___u4___fract_out_rnd2a;
	wire fpu___u4___exp_rnd_adj0;
	wire fpu___u4___exp_rnd_adj2a;
	wire fpu___u4___r_sign;
	wire fpu___u4___ovf0;
	wire fpu___u4___ovf1;
	wire [23:0] fpu___u4___fract_out_pl1;
	wire [7:0] fpu___u4___exp_out_pl1;
	wire [7:0] fpu___u4___exp_out_mi1;
	wire fpu___u4___exp_out_00;
	wire fpu___u4___exp_out_fe;
	wire fpu___u4___exp_out_ff;
	wire fpu___u4___exp_in_00;
	wire fpu___u4___exp_in_ff;
	wire fpu___u4___exp_out_final_ff;
	wire fpu___u4___fract_out_7fffff;
	wire [24:0] fpu___u4___fract_trunc;
	wire [7:0] fpu___u4___exp_out1;
	wire fpu___u4___grs_sel;
	wire fpu___u4___fract_out_00;
	wire fpu___u4___fract_in_00;
	wire fpu___u4___shft_co;
	wire [8:0] fpu___u4___exp_in_pl1;
	wire [8:0] fpu___u4___exp_in_mi1;
	wire [47:0] fpu___u4___fract_in_shftr;
	wire [47:0] fpu___u4___fract_in_shftl;
	wire [7:0] fpu___u4___exp_div;
	wire [7:0] fpu___u4___shft2;
	wire [7:0] fpu___u4___exp_out1_mi1;
	wire fpu___u4___div_dn;
	wire fpu___u4___div_nr;
	wire fpu___u4___grs_sel_div;
	wire fpu___u4___div_inf;
	wire [6:0] fpu___u4___fi_ldz_2a;
	wire [7:0] fpu___u4___fi_ldz_2;
	wire [7:0] fpu___u4___div_shft1;
	wire [7:0] fpu___u4___div_shft2;
	wire [7:0] fpu___u4___div_shft3;
	wire [7:0] fpu___u4___div_shft4;
	wire fpu___u4___div_shft1_co;
	wire [8:0] fpu___u4___div_exp1;
	wire [7:0] fpu___u4___div_exp2;
	wire [7:0] fpu___u4___div_exp3;
	wire fpu___u4___left_right;
	wire fpu___u4___lr_mul;
	wire fpu___u4___lr_div;
	wire [7:0] fpu___u4___shift_right;
	wire [7:0] fpu___u4___shftr_mul;
	wire [7:0] fpu___u4___shftr_div;
	wire [7:0] fpu___u4___shift_left;
	wire [7:0] fpu___u4___shftl_mul;
	wire [7:0] fpu___u4___shftl_div;
	wire [7:0] fpu___u4___fasu_shift;
	wire [7:0] fpu___u4___exp_fix_div;
	wire [7:0] fpu___u4___exp_fix_diva;
	wire [7:0] fpu___u4___exp_fix_divb;
	wire [5:0] fpu___u4___fi_ldz_mi1;
	wire [5:0] fpu___u4___fi_ldz_mi22;
	wire fpu___u4___exp_zero;
	wire [6:0] fpu___u4___ldz_all;
	wire [7:0] fpu___u4___ldz_dif;
	wire [8:0] fpu___u4___div_scht1a;
	wire [7:0] fpu___u4___f2i_shft;
	wire [55:0] fpu___u4___exp_f2i_1;
	wire fpu___u4___f2i_zero;
	wire fpu___u4___f2i_max;
	wire [7:0] fpu___u4___f2i_emin;
	wire [7:0] fpu___u4___conv_shft;
	wire [7:0] fpu___u4___exp_i2f;
	wire [7:0] fpu___u4___exp_f2i;
	wire [7:0] fpu___u4___conv_exp;
	wire fpu___u4___round2_f2i;
	wire fpu___u4___exp_in_80;
	wire fpu___u4___rmode_00;
	wire fpu___u4___rmode_01;
	wire fpu___u4___rmode_10;
	wire fpu___u4___rmode_11;
	parameter [7:0] fpu___u4___f2i_emax = 8'h9d;
	wire fpu___u4___max_num;
	wire fpu___u4___inf_out;
	wire fpu___u4___underflow_fmul;
	wire fpu___u4___overflow_fdiv;
	wire fpu___u4___undeflow_div;
	wire fpu___u4___z;
	wire fpu___u4___f2i_ine;
	assign fpu___clk = clk;
	assign fpu___rmode = rmode;
	assign fpu___fpu_op = fpu_op;
	assign fpu___opa = opa;
	assign fpu___opb = opb;
	assign fpu___sender_valid = sender_valid;
	wire [32:1] sv2v_tmp_CBA4B;
	assign sv2v_tmp_CBA4B = out;
	always @(*) fpu___out = sv2v_tmp_CBA4B;
	wire [1:1] sv2v_tmp_EDBAB;
	assign sv2v_tmp_EDBAB = inf;
	always @(*) fpu___inf = sv2v_tmp_EDBAB;
	wire [1:1] sv2v_tmp_5BCD5;
	assign sv2v_tmp_5BCD5 = snan;
	always @(*) fpu___snan = sv2v_tmp_5BCD5;
	wire [1:1] sv2v_tmp_AF4F5;
	assign sv2v_tmp_AF4F5 = qnan;
	always @(*) fpu___qnan = sv2v_tmp_AF4F5;
	wire [1:1] sv2v_tmp_A396B;
	assign sv2v_tmp_A396B = ine;
	always @(*) fpu___ine = sv2v_tmp_A396B;
	wire [1:1] sv2v_tmp_D5B3D;
	assign sv2v_tmp_D5B3D = overflow;
	always @(*) fpu___overflow = sv2v_tmp_D5B3D;
	wire [1:1] sv2v_tmp_1BC3F;
	assign sv2v_tmp_1BC3F = underflow;
	always @(*) fpu___underflow = sv2v_tmp_1BC3F;
	wire [1:1] sv2v_tmp_57FF5;
	assign sv2v_tmp_57FF5 = zero;
	always @(*) fpu___zero = sv2v_tmp_57FF5;
	wire [1:1] sv2v_tmp_AA3DB;
	assign sv2v_tmp_AA3DB = div_by_zero;
	always @(*) fpu___div_by_zero = sv2v_tmp_AA3DB;
	wire [1:1] sv2v_tmp_60C5B;
	assign sv2v_tmp_60C5B = input_ready;
	always @(*) fpu___input_ready = sv2v_tmp_60C5B;
	wire [1:1] sv2v_tmp_BA325;
	assign sv2v_tmp_BA325 = output_valid;
	always @(*) fpu___output_valid = sv2v_tmp_BA325;
	always @(posedge clk) begin
		input_ready <= 1'h1;
		fpu___data_accept_r1 <= input_ready & sender_valid;
		fpu___data_accept_r2 <= fpu___data_accept_r1;
		fpu___data_accept_r3 <= fpu___data_accept_r2;
		output_valid <= fpu___data_accept_r3;
	end
	always @(posedge clk) fpu___opa_r <= opa;
	always @(posedge clk) fpu___opb_r <= opb;
	always @(posedge clk) fpu___rmode_r1 <= rmode;
	always @(posedge clk) fpu___rmode_r2 <= fpu___rmode_r1;
	always @(posedge clk) fpu___rmode_r3 <= fpu___rmode_r2;
	always @(posedge clk) fpu___fpu_op_r1 <= fpu_op;
	always @(posedge clk) fpu___fpu_op_r2 <= fpu___fpu_op_r1;
	always @(posedge clk) fpu___fpu_op_r3 <= fpu___fpu_op_r2;
	assign fpu_____Vcellinp__u1__add = ~fpu___fpu_op_r1[2'h0+:32'h00000001];
	always @(posedge clk) fpu___sign_fasu_r <= fpu___sign_fasu;
	always @(posedge clk) fpu___sign_mul_r <= fpu___sign_mul;
	always @(posedge clk) fpu___sign_exe_r <= fpu___sign_exe;
	always @(posedge clk) fpu___inf_mul_r <= fpu___inf_mul;
	always @(posedge clk) fpu___exp_ovf_r <= fpu___exp_ovf;
	always @(posedge clk) fpu___fract_out_q <= {fpu___co_d, fpu___fract_out_d};
	always @(fpu___fracta_mul)
		case (fpu___fracta_mul[5'h00+:32'h00000017])
			23'b1zzzzzzzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h01;
			23'b01zzzzzzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h02;
			23'b001zzzzzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h03;
			23'b0001zzzzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h04;
			23'b00001zzzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h05;
			23'b000001zzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h06;
			23'b0000001zzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h07;
			23'b00000001zzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h08;
			23'b000000001zzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h09;
			23'b0000000001zzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h0a;
			23'b00000000001zzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h0b;
			23'b000000000001zzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h0c;
			23'b0000000000001zzzzzzzzzz: fpu___div_opa_ldz_d = 5'h0d;
			23'b00000000000001zzzzzzzzz: fpu___div_opa_ldz_d = 5'h0e;
			23'b000000000000001zzzzzzzz: fpu___div_opa_ldz_d = 5'h0f;
			23'b0000000000000001zzzzzzz: fpu___div_opa_ldz_d = 5'h10;
			23'b00000000000000001zzzzzz: fpu___div_opa_ldz_d = 5'h11;
			23'b000000000000000001zzzzz: fpu___div_opa_ldz_d = 5'h12;
			23'b0000000000000000001zzzz: fpu___div_opa_ldz_d = 5'h13;
			23'b00000000000000000001zzz: fpu___div_opa_ldz_d = 5'h14;
			23'b000000000000000000001zz: fpu___div_opa_ldz_d = 5'h15;
			23'b0000000000000000000001z: fpu___div_opa_ldz_d = 5'h16;
			23'bzzzzzzzzzzzzzzzzzzzzzzz: fpu___div_opa_ldz_d = 5'h17;
		endcase
	assign fpu___fdiv_opa = (|fpu___opa_r[5'h17+:32'h00000008] ? {fpu___fracta_mul, 26'h0000000} : {fpu___fracta_mul << fpu___div_opa_ldz_d, 26'h0000000});
	assign fpu___remainder = {26'b00000000000000000000000000, fpu_____Vcellout__u_divider__remainder};
	assign fpu___remainder_00 = ~(|fpu___remainder);
	always @(posedge clk) fpu___div_opa_ldz_r1 <= fpu___div_opa_ldz_d;
	always @(posedge clk) fpu___div_opa_ldz_r2 <= fpu___div_opa_ldz_r1;
	always @(posedge clk)
		case ({29'b00000000000000000000000000000, fpu___fpu_op_r2})
			32'sh00000000, 32'sh00000001: fpu___exp_r <= fpu___exp_fasu;
			32'sh00000002, 32'sh00000003: fpu___exp_r <= fpu___exp_mul;
			32'sh00000004: fpu___exp_r <= 8'h00;
			32'sh00000005: fpu___exp_r <= fpu___opa_r1[5'h17+:32'h00000008];
		endcase
	assign fpu___fract_div = (fpu___opb_dn ? fpu___quo[6'h02+:32'h00000030] : {fpu___quo[6'h00+:32'h0000001b], 21'h000000});
	always @(posedge clk) fpu___opa_r1 <= fpu___opa_r[5'h00+:32'h0000001f];
	always @(posedge clk) fpu___fract_i2f <= (3'h5 == fpu___fpu_op_r2 ? (fpu___sign_d ? (48'h000000000001 - {24'b000000000000000000000000, |fpu___opa_r1[5'h17+:32'h00000008], fpu___opa_r1[5'h00+:32'h00000017]}) - 48'h000000000001 : {24'b000000000000000000000000, |fpu___opa_r1[5'h17+:32'h00000008], fpu___opa_r1[5'h00+:32'h00000017]}) : (fpu___sign_d ? 48'h000000000001 - {fpu___opa_r1, 17'h00001} : {fpu___opa_r1, 17'h00000}));
	always @(fpu___fpu_op_r3 or fpu___fract_div or fpu___fract_i2f or fpu___fract_out_q or fpu___prod)
		case ({29'b00000000000000000000000000000, fpu___fpu_op_r3})
			32'sh00000000, 32'sh00000001: fpu___fract_denorm = {fpu___fract_out_q, 20'h00000};
			32'sh00000002: fpu___fract_denorm = fpu___prod;
			32'sh00000003: fpu___fract_denorm = fpu___fract_div;
			32'sh00000004, 32'sh00000005: fpu___fract_denorm = fpu___fract_i2f;
			default: fpu___fract_denorm = 48'h000000000000;
		endcase
	always @(posedge clk) fpu___opas_r1 <= fpu___opa_r[5'h1f+:32'h00000001];
	always @(posedge clk) fpu___opas_r2 <= fpu___opas_r1;
	assign fpu___sign_d = (fpu___fpu_op_r2[2'h1+:32'h00000001] ? fpu___sign_mul : fpu___sign_fasu);
	always @(posedge clk) fpu___sign <= (2'h3 == fpu___rmode_r2 ? ~fpu___sign_d : fpu___sign_d);
	assign fpu_____Vcellinp__u4__output_zero = fpu___mul_00 | fpu___div_00;
	always @(posedge clk) fpu___fasu_op_r1 <= fpu___fasu_op;
	always @(posedge clk) fpu___fasu_op_r2 <= fpu___fasu_op_r1;
	always @(posedge clk) fpu___inf_mul2 <= 8'hff == fpu___exp_mul;
	assign fpu___mul_inf = ((3'h2 == fpu___fpu_op_r3) & (fpu___inf_mul_r | fpu___inf_mul2)) & (2'h0 == fpu___rmode_r3);
	assign fpu___div_inf = (3'h3 == fpu___fpu_op_r3) & (fpu___opb_00 | fpu___opa_inf);
	assign fpu___mul_00 = (3'h2 == fpu___fpu_op_r3) & (fpu___opa_00 | fpu___opb_00);
	assign fpu___div_00 = (3'h3 == fpu___fpu_op_r3) & (fpu___opa_00 | fpu___opb_inf);
	assign fpu___out_fixed = ((((fpu___qnan_d | fpu___snan_d) | (fpu___ind_d & ~fpu___fasu_op_r2)) | (((3'h3 == fpu___fpu_op_r3) & fpu___opb_00) & fpu___opa_00)) | (((fpu___opa_inf & fpu___opb_00) | (fpu___opb_inf & fpu___opa_00)) & (3'h2 == fpu___fpu_op_r3)) ? 31'h7fc00001 : 31'h7f800000);
	always @(posedge clk) out[5'h00+:32'h0000001f] <= (((((fpu___mul_inf | fpu___div_inf) | ((fpu___inf_d & (3'h3 != fpu___fpu_op_r3)) & (3'h5 != fpu___fpu_op_r3))) | fpu___snan_d) | fpu___qnan_d) & (3'h4 != fpu___fpu_op_r3) ? fpu___out_fixed : fpu___out_d);
	assign fpu___out_d_00 = ~(|fpu___out_d);
	assign fpu___sign_mul_final = (fpu___sign_exe_r & ((fpu___opa_00 & fpu___opb_inf) | (fpu___opb_00 & fpu___opa_inf)) ? ~fpu___sign_mul_r : fpu___sign_mul_r);
	assign fpu___sign_div_final = (fpu___sign_exe_r & (fpu___opa_inf & fpu___opb_inf) ? ~fpu___sign_mul_r : fpu___sign_mul_r | (fpu___opa_00 & fpu___opb_00));
	always @(posedge clk) out[5'h1f+:32'h00000001] <= ((3'h5 == fpu___fpu_op_r3) & fpu___out_d_00 ? fpu___f2i_out_sign & ~(fpu___qnan_d | fpu___snan_d) : ((3'h2 == fpu___fpu_op_r3) & ~(fpu___snan_d | fpu___qnan_d) ? fpu___sign_mul_final : ((3'h3 == fpu___fpu_op_r3) & ~(fpu___snan_d | fpu___qnan_d) ? fpu___sign_div_final : ((fpu___snan_d | fpu___qnan_d) | fpu___ind_d ? fpu___nan_sign_d : (fpu___output_zero_fasu ? fpu___result_zero_sign_d : fpu___sign_fasu_r)))));
	assign fpu___ine_mula = (((((fpu___inf_mul_r | fpu___inf_mul2) | fpu___opa_inf) | fpu___opb_inf) & (2'h1 == fpu___rmode_r3)) & ~((fpu___opa_inf & fpu___opb_00) | (fpu___opb_inf & fpu___opa_00))) & fpu___fpu_op_r3[2'h1+:32'h00000001];
	assign fpu___ine_mul = (((((((fpu___ine_mula | fpu___ine_d) | fpu___inf_fmul) | fpu___out_d_00) | fpu___overflow_d) | fpu___underflow_d) & ~fpu___opa_00) & ~fpu___opb_00) & ~((fpu___snan_d | fpu___qnan_d) | fpu___inf_d);
	assign fpu___ine_div = ((fpu___ine_d | fpu___overflow_d) | fpu___underflow_d) & ~(((fpu___opb_00 | fpu___snan_d) | fpu___qnan_d) | fpu___inf_d);
	assign fpu___ine_fasu = ((fpu___ine_d | fpu___overflow_d) | fpu___underflow_d) & ~((fpu___snan_d | fpu___qnan_d) | fpu___inf_d);
	always @(posedge clk) ine <= (fpu___fpu_op_r3[2'h2+:32'h00000001] ? fpu___ine_d : (fpu___fpu_op_r3[2'h1+:32'h00000001] ? (fpu___fpu_op_r3[2'h0+:32'h00000001] ? fpu___ine_div : fpu___ine_mul) : fpu___ine_fasu));
	assign fpu___overflow_fasu = fpu___overflow_d & ~((fpu___snan_d | fpu___qnan_d) | fpu___inf_d);
	assign fpu___overflow_fmul = (~fpu___inf_d & ((fpu___inf_mul_r | fpu___inf_mul2) | fpu___overflow_d)) & ~(fpu___snan_d | fpu___qnan_d);
	assign fpu___overflow_fdiv = fpu___overflow_d & ~(((fpu___opb_00 | fpu___inf_d) | fpu___snan_d) | fpu___qnan_d);
	always @(posedge clk) begin
		___sel_temp_0 = (fpu___fpu_op_r3[2'h2+:32'h00000001] ? 32'sh00000000 : (fpu___fpu_op_r3[2'h1+:32'h00000001] ? (fpu___fpu_op_r3[2'h0+:32'h00000001] ? {31'b0000000000000000000000000000000, fpu___overflow_fdiv} : {31'b0000000000000000000000000000000, fpu___overflow_fmul}) : {31'b0000000000000000000000000000000, fpu___overflow_fasu}));
		overflow <= ___sel_temp_0[32'h00000000+:32'h00000001];
	end
	always @(posedge clk) fpu___underflow_fmul_r <= fpu___underflow_fmul_d;
	assign fpu___underflow_fmul1 = ((fpu___underflow_fmul_r[2'h0+:32'h00000001] | (fpu___underflow_fmul_r[2'h1+:32'h00000001] & fpu___underflow_d)) | ((((fpu___opa_dn | fpu___opb_dn) & fpu___out_d_00) & (48'h000000000000 != fpu___prod)) & fpu___sign)) | (fpu___underflow_fmul_r[2'h2+:32'h00000001] & ((8'h00 == fpu___out_d[5'h17+:32'h00000008]) | (23'h000000 == fpu___out_d[5'h00+:32'h00000017])));
	assign fpu___underflow_fasu = fpu___underflow_d & ~((fpu___inf_d | fpu___snan_d) | fpu___qnan_d);
	assign fpu___underflow_fmul = fpu___underflow_fmul1 & ~((fpu___snan_d | fpu___qnan_d) | fpu___inf_mul_r);
	assign fpu___underflow_fdiv = fpu___underflow_fasu & ~fpu___opb_00;
	always @(posedge clk) begin
		___sel_temp_1 = (fpu___fpu_op_r3[2'h2+:32'h00000001] ? 32'sh00000000 : (fpu___fpu_op_r3[2'h1+:32'h00000001] ? (fpu___fpu_op_r3[2'h0+:32'h00000001] ? {31'b0000000000000000000000000000000, fpu___underflow_fdiv} : {31'b0000000000000000000000000000000, fpu___underflow_fmul}) : {31'b0000000000000000000000000000000, fpu___underflow_fasu}));
		underflow <= ___sel_temp_1[32'h00000000+:32'h00000001];
	end
	always @(posedge clk) snan <= fpu___snan_d;
	always @(posedge clk) begin
		___sel_temp_2 = (fpu___fpu_op_r3[2'h2+:32'h00000001] ? 32'sh00000000 : ((({31'b0000000000000000000000000000000, fpu___snan_d} | {31'b0000000000000000000000000000000, fpu___qnan_d}) | ({31'b0000000000000000000000000000000, fpu___ind_d} & {31'b0000000000000000000000000000000, ~fpu___fasu_op_r2})) | (({31'b0000000000000000000000000000000, fpu___opa_00} & {31'b0000000000000000000000000000000, fpu___opb_00}) & {31'b0000000000000000000000000000000, 3'h3 == fpu___fpu_op_r3})) | ((({31'b0000000000000000000000000000000, fpu___opa_inf} & {31'b0000000000000000000000000000000, fpu___opb_00}) | ({31'b0000000000000000000000000000000, fpu___opb_inf} & {31'b0000000000000000000000000000000, fpu___opa_00})) & {31'b0000000000000000000000000000000, 3'h2 == fpu___fpu_op_r3}));
		qnan <= ___sel_temp_2[32'h00000000+:32'h00000001];
	end
	assign fpu___inf_fmul = (((((fpu___inf_mul_r | fpu___inf_mul2) & (2'h0 == fpu___rmode_r3)) | fpu___opa_inf) | fpu___opb_inf) & ~((fpu___opa_inf & fpu___opb_00) | (fpu___opb_inf & fpu___opa_00))) & (3'h2 == fpu___fpu_op_r3);
	always @(posedge clk) begin
		___sel_temp_3 = (fpu___fpu_op_r3[2'h2+:32'h00000001] ? 32'sh00000000 : {31'b0000000000000000000000000000000, ~(fpu___qnan_d | fpu___snan_d)} & (((((({31'b0000000000000000000000000000000, &fpu___out_d[5'h17+:32'h00000008]} & {31'b0000000000000000000000000000000, ~(|fpu___out_d[5'h00+:32'h00000017])}) & {31'b0000000000000000000000000000000, ~(fpu___opb_00 & (3'h3 == fpu___fpu_op_r3))}) | (({31'b0000000000000000000000000000000, fpu___inf_d} & {31'b0000000000000000000000000000000, ~(fpu___ind_d & ~fpu___fasu_op_r2)}) & {31'b0000000000000000000000000000000, ~fpu___fpu_op_r3[2'h1+:32'h00000001]})) | {31'b0000000000000000000000000000000, fpu___inf_fmul}) | (({31'b0000000000000000000000000000000, ~fpu___opa_00} & {31'b0000000000000000000000000000000, fpu___opb_00}) & {31'b0000000000000000000000000000000, 3'h3 == fpu___fpu_op_r3})) | (({31'b0000000000000000000000000000000, 3'h3 == fpu___fpu_op_r3} & {31'b0000000000000000000000000000000, fpu___opa_inf}) & {31'b0000000000000000000000000000000, ~fpu___opb_inf})));
		inf <= ___sel_temp_3[32'h00000000+:32'h00000001];
	end
	assign fpu___output_zero_fasu = fpu___out_d_00 & ~((fpu___inf_d | fpu___snan_d) | fpu___qnan_d);
	assign fpu___output_zero_fdiv = (((fpu___div_00 | (fpu___out_d_00 & ~fpu___opb_00)) & ~(fpu___opa_inf & fpu___opb_inf)) & ~(fpu___opa_00 & fpu___opb_00)) & ~(fpu___qnan_d | fpu___snan_d);
	assign fpu___output_zero_fmul = ((((fpu___out_d_00 | fpu___opa_00) | fpu___opb_00) & ~(((((fpu___inf_mul_r | fpu___inf_mul2) | fpu___opa_inf) | fpu___opb_inf) | fpu___snan_d) | fpu___qnan_d)) & ~(fpu___opa_inf & fpu___opb_00)) & ~(fpu___opb_inf & fpu___opa_00);
	always @(posedge clk) zero <= (3'h5 == fpu___fpu_op_r3 ? fpu___out_d_00 & ~(fpu___snan_d | fpu___qnan_d) : (3'h3 == fpu___fpu_op_r3 ? fpu___output_zero_fdiv : (3'h2 == fpu___fpu_op_r3 ? fpu___output_zero_fmul : fpu___output_zero_fasu)));
	always @(posedge clk) fpu___opa_nan_r <= ~fpu___opa_nan & (3'h3 == fpu___fpu_op_r2);
	always @(posedge clk) div_by_zero <= ((fpu___opa_nan_r & ~fpu___opa_00) & ~fpu___opa_inf) & fpu___opb_00;
	assign fpu___u0___clk = fpu___clk;
	assign fpu___u0___opa = fpu___opa_r;
	assign fpu___u0___opb = fpu___opb_r;
	wire [1:1] sv2v_tmp_761B5;
	assign sv2v_tmp_761B5 = fpu___inf_d;
	always @(*) fpu___u0___inf = sv2v_tmp_761B5;
	wire [1:1] sv2v_tmp_60175;
	assign sv2v_tmp_60175 = fpu___ind_d;
	always @(*) fpu___u0___ind = sv2v_tmp_60175;
	wire [1:1] sv2v_tmp_48D57;
	assign sv2v_tmp_48D57 = fpu___qnan_d;
	always @(*) fpu___u0___qnan = sv2v_tmp_48D57;
	wire [1:1] sv2v_tmp_F9CF7;
	assign sv2v_tmp_F9CF7 = fpu___snan_d;
	always @(*) fpu___u0___snan = sv2v_tmp_F9CF7;
	wire [1:1] sv2v_tmp_69520;
	assign sv2v_tmp_69520 = fpu___opa_nan;
	always @(*) fpu___u0___opa_nan = sv2v_tmp_69520;
	wire [1:1] sv2v_tmp_E10A0;
	assign sv2v_tmp_E10A0 = fpu___opb_nan;
	always @(*) fpu___u0___opb_nan = sv2v_tmp_E10A0;
	wire [1:1] sv2v_tmp_E54D2;
	assign sv2v_tmp_E54D2 = fpu___opa_00;
	always @(*) fpu___u0___opa_00 = sv2v_tmp_E54D2;
	wire [1:1] sv2v_tmp_04582;
	assign sv2v_tmp_04582 = fpu___opb_00;
	always @(*) fpu___u0___opb_00 = sv2v_tmp_04582;
	wire [1:1] sv2v_tmp_79BE0;
	assign sv2v_tmp_79BE0 = fpu___opa_inf;
	always @(*) fpu___u0___opa_inf = sv2v_tmp_79BE0;
	wire [1:1] sv2v_tmp_72A80;
	assign sv2v_tmp_72A80 = fpu___opb_inf;
	always @(*) fpu___u0___opb_inf = sv2v_tmp_72A80;
	wire [1:1] sv2v_tmp_50252;
	assign sv2v_tmp_50252 = fpu___opa_dn;
	always @(*) fpu___u0___opa_dn = sv2v_tmp_50252;
	wire [1:1] sv2v_tmp_51962;
	assign sv2v_tmp_51962 = fpu___opb_dn;
	always @(*) fpu___u0___opb_dn = sv2v_tmp_51962;
	assign fpu___u0___expa = fpu___opa_r[5'h17+:32'h00000008];
	assign fpu___u0___expb = fpu___opb_r[5'h17+:32'h00000008];
	assign fpu___u0___fracta = fpu___opa_r[5'h00+:32'h00000017];
	assign fpu___u0___fractb = fpu___opb_r[5'h00+:32'h00000017];
	always @(posedge clk) fpu___u0___expa_ff <= &fpu___u0___expa;
	always @(posedge clk) fpu___u0___expb_ff <= &fpu___u0___expb;
	always @(posedge clk) fpu___u0___infa_f_r <= ~(|fpu___u0___fracta);
	always @(posedge clk) fpu___u0___infb_f_r <= ~(|fpu___u0___fractb);
	always @(posedge clk) fpu___u0___qnan_r_a <= fpu___u0___fracta[5'h16+:32'h00000001];
	always @(posedge clk) fpu___u0___snan_r_a <= ~fpu___u0___fracta[5'h16+:32'h00000001] & |fpu___u0___fracta[5'h00+:32'h00000016];
	always @(posedge clk) fpu___u0___qnan_r_b <= fpu___u0___fractb[5'h16+:32'h00000001];
	always @(posedge clk) fpu___u0___snan_r_b <= ~fpu___u0___fractb[5'h16+:32'h00000001] & |fpu___u0___fractb[5'h00+:32'h00000016];
	always @(posedge clk) fpu___ind_d <= (fpu___u0___expa_ff & fpu___u0___infa_f_r) & (fpu___u0___expb_ff & fpu___u0___infb_f_r);
	always @(posedge clk) fpu___inf_d <= (fpu___u0___expa_ff & fpu___u0___infa_f_r) | (fpu___u0___expb_ff & fpu___u0___infb_f_r);
	always @(posedge clk) fpu___qnan_d <= (fpu___u0___expa_ff & fpu___u0___qnan_r_a) | (fpu___u0___expb_ff & fpu___u0___qnan_r_b);
	always @(posedge clk) fpu___snan_d <= (fpu___u0___expa_ff & fpu___u0___snan_r_a) | (fpu___u0___expb_ff & fpu___u0___snan_r_b);
	always @(posedge clk) fpu___opa_nan <= &fpu___u0___expa & |fpu___u0___fracta;
	always @(posedge clk) fpu___opb_nan <= &fpu___u0___expb & |fpu___u0___fractb;
	always @(posedge clk) fpu___opa_inf <= fpu___u0___expa_ff & fpu___u0___infa_f_r;
	always @(posedge clk) fpu___opb_inf <= fpu___u0___expb_ff & fpu___u0___infb_f_r;
	always @(posedge clk) fpu___u0___expa_00 <= ~(|fpu___u0___expa);
	always @(posedge clk) fpu___u0___expb_00 <= ~(|fpu___u0___expb);
	always @(posedge clk) fpu___u0___fracta_00 <= ~(|fpu___u0___fracta);
	always @(posedge clk) fpu___u0___fractb_00 <= ~(|fpu___u0___fractb);
	always @(posedge clk) fpu___opa_00 <= fpu___u0___expa_00 & fpu___u0___fracta_00;
	always @(posedge clk) fpu___opb_00 <= fpu___u0___expb_00 & fpu___u0___fractb_00;
	always @(posedge clk) fpu___opa_dn <= fpu___u0___expa_00;
	always @(posedge clk) fpu___opb_dn <= fpu___u0___expb_00;
	assign fpu___u1___clk = fpu___clk;
	assign fpu___u1___rmode = fpu___rmode_r2;
	assign fpu___u1___add = fpu_____Vcellinp__u1__add;
	assign fpu___u1___opa = fpu___opa_r;
	assign fpu___u1___opb = fpu___opb_r;
	assign fpu___u1___opa_nan = fpu___opa_nan;
	assign fpu___u1___opb_nan = fpu___opb_nan;
	wire [27:1] sv2v_tmp_28A36;
	assign sv2v_tmp_28A36 = fpu___fracta;
	always @(*) fpu___u1___fracta_out = sv2v_tmp_28A36;
	wire [27:1] sv2v_tmp_F2CC6;
	assign sv2v_tmp_F2CC6 = fpu___fractb;
	always @(*) fpu___u1___fractb_out = sv2v_tmp_F2CC6;
	wire [8:1] sv2v_tmp_1853F;
	assign sv2v_tmp_1853F = fpu___exp_fasu;
	always @(*) fpu___u1___exp_dn_out = sv2v_tmp_1853F;
	wire [1:1] sv2v_tmp_0C0FC;
	assign sv2v_tmp_0C0FC = fpu___sign_fasu;
	always @(*) fpu___u1___sign = sv2v_tmp_0C0FC;
	wire [1:1] sv2v_tmp_1539E;
	assign sv2v_tmp_1539E = fpu___nan_sign_d;
	always @(*) fpu___u1___nan_sign = sv2v_tmp_1539E;
	wire [1:1] sv2v_tmp_A5EDE;
	assign sv2v_tmp_A5EDE = fpu___result_zero_sign_d;
	always @(*) fpu___u1___result_zero_sign = sv2v_tmp_A5EDE;
	wire [1:1] sv2v_tmp_76201;
	assign sv2v_tmp_76201 = fpu___fasu_op;
	always @(*) fpu___u1___fasu_op = sv2v_tmp_76201;
	assign fpu___u1___signa = fpu___opa_r[5'h1f+:32'h00000001];
	assign fpu___u1___signb = fpu___opb_r[5'h1f+:32'h00000001];
	assign fpu___u1___expa = fpu___opa_r[5'h17+:32'h00000008];
	assign fpu___u1___expb = fpu___opb_r[5'h17+:32'h00000008];
	assign fpu___u1___fracta = fpu___opa_r[5'h00+:32'h00000017];
	assign fpu___u1___fractb = fpu___opb_r[5'h00+:32'h00000017];
	assign fpu___u1___expa_lt_expb = fpu___u1___expa > fpu___u1___expb;
	assign fpu___u1___expa_dn = ~(|fpu___u1___expa);
	assign fpu___u1___expb_dn = ~(|fpu___u1___expb);
	assign fpu___u1___exp_small = (fpu___u1___expa_lt_expb ? fpu___u1___expb : fpu___u1___expa);
	assign fpu___u1___exp_large = (fpu___u1___expa_lt_expb ? fpu___u1___expa : fpu___u1___expb);
	assign fpu___u1___exp_diff1 = fpu___u1___exp_large - fpu___u1___exp_small;
	assign fpu___u1___exp_diff1a = fpu___u1___exp_diff1 - 8'h01;
	assign fpu___u1___exp_diff2 = (fpu___u1___expa_dn | fpu___u1___expb_dn ? fpu___u1___exp_diff1a : fpu___u1___exp_diff1);
	assign fpu___u1___exp_diff = (fpu___u1___expa_dn & fpu___u1___expb_dn ? 8'h00 : fpu___u1___exp_diff2);
	always @(posedge clk) fpu___exp_fasu <= ((~fpu___u1___add_d & (fpu___u1___expa == fpu___u1___expb)) & (fpu___u1___fracta == fpu___u1___fractb) ? 8'h00 : fpu___u1___exp_large);
	assign fpu___u1___op_dn = (fpu___u1___expa_lt_expb ? fpu___u1___expb_dn : fpu___u1___expa_dn);
	assign fpu___u1___adj_op = (fpu___u1___expa_lt_expb ? fpu___u1___fractb : fpu___u1___fracta);
	assign fpu___u1___adj_op_tmp = {~fpu___u1___op_dn, fpu___u1___adj_op, 3'h0};
	assign fpu___u1___exp_lt_27 = 8'h1b < fpu___u1___exp_diff;
	assign fpu___u1___exp_diff_sft = (fpu___u1___exp_lt_27 ? 5'h1b : fpu___u1___exp_diff[3'h0+:32'h00000005]);
	assign fpu___u1___adj_op_out_sft = fpu___u1___adj_op_tmp >> fpu___u1___exp_diff_sft;
	assign fpu___u1___adj_op_out = {fpu___u1___adj_op_out_sft[5'h01+:32'h0000001a], fpu___u1___adj_op_out_sft[5'h00+:32'h00000001] | fpu___u1___sticky};
	always @(fpu___u1___adj_op_tmp or fpu___u1___exp_diff_sft)
		case ({27'b000000000000000000000000000, fpu___u1___exp_diff_sft})
			32'sh00000000: fpu___u1___sticky = 1'h0;
			32'sh00000001: fpu___u1___sticky = fpu___u1___adj_op_tmp[5'h00+:32'h00000001];
			32'sh00000002: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000002];
			32'sh00000003: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000003];
			32'sh00000004: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000004];
			32'sh00000005: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000005];
			32'sh00000006: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000006];
			32'sh00000007: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000007];
			32'sh00000008: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000008];
			32'sh00000009: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000009];
			32'sh0000000a: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000000a];
			32'sh0000000b: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000000b];
			32'sh0000000c: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000000c];
			32'sh0000000d: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000000d];
			32'sh0000000e: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000000e];
			32'sh0000000f: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000000f];
			32'sh00000010: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000010];
			32'sh00000011: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000011];
			32'sh00000012: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000012];
			32'sh00000013: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000013];
			32'sh00000014: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000014];
			32'sh00000015: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000015];
			32'sh00000016: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000016];
			32'sh00000017: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000017];
			32'sh00000018: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000018];
			32'sh00000019: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h00000019];
			32'sh0000001a: fpu___u1___sticky = |fpu___u1___adj_op_tmp[5'h00+:32'h0000001a];
			32'sh0000001b: fpu___u1___sticky = |fpu___u1___adj_op_tmp;
		endcase
	assign fpu___u1___fracta_n = (fpu___u1___expa_lt_expb ? {~fpu___u1___expa_dn, fpu___u1___fracta, 3'h0} : fpu___u1___adj_op_out);
	assign fpu___u1___fractb_n = (fpu___u1___expa_lt_expb ? fpu___u1___adj_op_out : {~fpu___u1___expb_dn, fpu___u1___fractb, 3'h0});
	assign fpu___u1___fractb_lt_fracta = fpu___u1___fractb_n > fpu___u1___fracta_n;
	assign fpu___u1___fracta_s = (fpu___u1___fractb_lt_fracta ? fpu___u1___fractb_n : fpu___u1___fracta_n);
	assign fpu___u1___fractb_s = (fpu___u1___fractb_lt_fracta ? fpu___u1___fracta_n : fpu___u1___fractb_n);
	always @(posedge clk) fpu___fracta <= fpu___u1___fracta_s;
	always @(posedge clk) fpu___fractb <= fpu___u1___fractb_s;
	always @(fpu_____Vcellinp__u1__add or fpu___u1___fractb_lt_fracta or fpu___u1___signa or fpu___u1___signb)
		case ({fpu___u1___signa, fpu___u1___signb, fpu_____Vcellinp__u1__add})
			3'h1: fpu___u1___sign_d = 1'h0;
			3'h3: fpu___u1___sign_d = fpu___u1___fractb_lt_fracta;
			3'h5: fpu___u1___sign_d = ~fpu___u1___fractb_lt_fracta;
			3'h7: fpu___u1___sign_d = 1'h1;
			3'h0: fpu___u1___sign_d = fpu___u1___fractb_lt_fracta;
			3'h2: fpu___u1___sign_d = 1'h0;
			3'h4: fpu___u1___sign_d = 1'h1;
			3'h6: fpu___u1___sign_d = ~fpu___u1___fractb_lt_fracta;
		endcase
	always @(posedge clk) fpu___sign_fasu <= fpu___u1___sign_d;
	always @(posedge clk) fpu___u1___signa_r <= fpu___u1___signa;
	always @(posedge clk) fpu___u1___signb_r <= fpu___u1___signb;
	always @(posedge clk) fpu___u1___add_r <= fpu_____Vcellinp__u1__add;
	always @(posedge clk) fpu___result_zero_sign_d <= ((((fpu___u1___add_r & fpu___u1___signa_r) & fpu___u1___signb_r) | ((~fpu___u1___add_r & fpu___u1___signa_r) & ~fpu___u1___signb_r)) | ((fpu___u1___add_r & (fpu___u1___signa_r | fpu___u1___signb_r)) & (2'h3 == fpu___rmode_r2))) | ((~fpu___u1___add_r & (fpu___u1___signa_r == fpu___u1___signb_r)) & (2'h3 == fpu___rmode_r2));
	always @(posedge clk) fpu___u1___fracta_lt_fractb <= fpu___u1___fracta < fpu___u1___fractb;
	always @(posedge clk) fpu___u1___fracta_eq_fractb <= fpu___u1___fracta == fpu___u1___fractb;
	assign fpu___u1___nan_sign1 = (fpu___u1___fracta_eq_fractb ? fpu___u1___signa_r & fpu___u1___signb_r : (fpu___u1___fracta_lt_fractb ? fpu___u1___signb_r : fpu___u1___signa_r));
	always @(posedge clk) fpu___nan_sign_d <= (fpu___opa_nan & fpu___opb_nan ? fpu___u1___nan_sign1 : (fpu___opb_nan ? fpu___u1___signb_r : fpu___u1___signa_r));
	always @(fpu_____Vcellinp__u1__add or fpu___u1___signa or fpu___u1___signb)
		case ({fpu___u1___signa, fpu___u1___signb, fpu_____Vcellinp__u1__add})
			3'h1: fpu___u1___add_d = 1'h1;
			3'h3: fpu___u1___add_d = 1'h0;
			3'h5: fpu___u1___add_d = 1'h0;
			3'h7: fpu___u1___add_d = 1'h1;
			3'h0: fpu___u1___add_d = 1'h0;
			3'h2: fpu___u1___add_d = 1'h1;
			3'h4: fpu___u1___add_d = 1'h1;
			3'h6: fpu___u1___add_d = 1'h0;
		endcase
	always @(posedge clk) fpu___fasu_op <= fpu___u1___add_d;
	assign fpu___u2___clk = fpu___clk;
	assign fpu___u2___fpu_op = fpu___fpu_op_r1;
	assign fpu___u2___opa = fpu___opa_r;
	assign fpu___u2___opb = fpu___opb_r;
	assign fpu___u2___fracta = fpu___fracta_mul;
	assign fpu___u2___fractb = fpu___fractb_mul;
	wire [8:1] sv2v_tmp_AF418;
	assign sv2v_tmp_AF418 = fpu___exp_mul;
	always @(*) fpu___u2___exp_out = sv2v_tmp_AF418;
	wire [1:1] sv2v_tmp_72C1B;
	assign sv2v_tmp_72C1B = fpu___sign_mul;
	always @(*) fpu___u2___sign = sv2v_tmp_72C1B;
	wire [1:1] sv2v_tmp_A2CA4;
	assign sv2v_tmp_A2CA4 = fpu___sign_exe;
	always @(*) fpu___u2___sign_exe = sv2v_tmp_A2CA4;
	wire [1:1] sv2v_tmp_A8F55;
	assign sv2v_tmp_A8F55 = fpu___inf_mul;
	always @(*) fpu___u2___inf = sv2v_tmp_A8F55;
	wire [2:1] sv2v_tmp_35DA2;
	assign sv2v_tmp_35DA2 = fpu___exp_ovf;
	always @(*) fpu___u2___exp_ovf = sv2v_tmp_35DA2;
	wire [3:1] sv2v_tmp_C3DCB;
	assign sv2v_tmp_C3DCB = fpu___underflow_fmul_d;
	always @(*) fpu___u2___underflow = sv2v_tmp_C3DCB;
	assign fpu___u2___op_div = 3'h3 == fpu___fpu_op_r1;
	assign fpu___u2___signa = fpu___opa_r[5'h1f+:32'h00000001];
	assign fpu___u2___signb = fpu___opb_r[5'h1f+:32'h00000001];
	assign fpu___u2___expa = fpu___opa_r[5'h17+:32'h00000008];
	assign fpu___u2___expb = fpu___opb_r[5'h17+:32'h00000008];
	assign fpu___u2___expa_dn = ~(|fpu___u2___expa);
	assign fpu___u2___expb_dn = ~(|fpu___u2___expb);
	assign fpu___u2___opa_00 = ~(|fpu___opa_r[5'h00+:32'h0000001f]);
	assign fpu___u2___opb_00 = ~(|fpu___opb_r[5'h00+:32'h0000001f]);
	assign fpu___u2___fracta_00 = ~(|fpu___opa_r[5'h00+:32'h00000017]);
	assign fpu___u2___fractb_00 = ~(|fpu___opb_r[5'h00+:32'h00000017]);
	assign fpu___fracta_mul = {~fpu___u2___expa_dn, fpu___opa_r[5'h00+:32'h00000017]};
	assign fpu___fractb_mul = {~fpu___u2___expb_dn, fpu___opb_r[5'h00+:32'h00000017]};
	assign ___sel_temp_4 = (fpu___u2___op_div ? {1'b0, fpu___u2___expa} - {1'b0, fpu___u2___expb} : {1'b0, fpu___u2___expa} + {1'b0, fpu___u2___expb});
	assign fpu___u2___co1 = ___sel_temp_4[32'h00000008+:32'h00000001];
	assign ___sel_temp_5 = (fpu___u2___op_div ? {1'b0, fpu___u2___expa} - {1'b0, fpu___u2___expb} : {1'b0, fpu___u2___expa} + {1'b0, fpu___u2___expb});
	assign fpu___u2___exp_tmp1 = ___sel_temp_5[32'h00000000+:32'h00000008];
	assign ___sel_temp_6 = (fpu___u2___op_div ? 9'h07f + {fpu___u2___co1, fpu___u2___exp_tmp1} : {fpu___u2___co1, fpu___u2___exp_tmp1} - 9'h07f);
	assign fpu___u2___co2 = ___sel_temp_6[32'h00000008+:32'h00000001];
	assign ___sel_temp_7 = (fpu___u2___op_div ? 9'h07f + {fpu___u2___co1, fpu___u2___exp_tmp1} : {fpu___u2___co1, fpu___u2___exp_tmp1} - 9'h07f);
	assign fpu___u2___exp_tmp2 = ___sel_temp_7[32'h00000000+:32'h00000008];
	assign fpu___u2___exp_tmp3 = 8'h01 + fpu___u2___exp_tmp2;
	assign fpu___u2___exp_tmp4 = 8'h7f - fpu___u2___exp_tmp1;
	assign ___sel_temp_8 = (fpu___u2___op_div ? 32'sh00000001 + {24'b000000000000000000000000, fpu___u2___exp_tmp4} : {24'b000000000000000000000000, fpu___u2___exp_tmp4} - 32'sh00000001);
	assign fpu___u2___exp_tmp5 = ___sel_temp_8[32'h00000000+:32'h00000008];
	always @(posedge clk) fpu___exp_mul <= (fpu___u2___op_div ? fpu___u2___exp_out_div : fpu___u2___exp_out_mul);
	assign fpu___u2___exp_out_div = (fpu___u2___expa_dn | fpu___u2___expb_dn ? (fpu___u2___co2 ? fpu___u2___exp_tmp5 : fpu___u2___exp_tmp3) : (fpu___u2___co2 ? fpu___u2___exp_tmp4 : fpu___u2___exp_tmp2));
	assign fpu___u2___exp_out_mul = (fpu___u2___exp_ovf_d[1'h1+:32'h00000001] ? fpu___u2___exp_out_a : (fpu___u2___expa_dn | fpu___u2___expb_dn ? fpu___u2___exp_tmp3 : fpu___u2___exp_tmp2));
	assign fpu___u2___exp_out_a = (fpu___u2___expa_dn | fpu___u2___expb_dn ? fpu___u2___exp_tmp5 : fpu___u2___exp_tmp4);
	assign fpu___u2___exp_ovf_d[1'h0+:32'h00000001] = (fpu___u2___op_div ? fpu___u2___expa[3'h7+:32'h00000001] & ~fpu___u2___expb[3'h7+:32'h00000001] : (fpu___u2___co2 & fpu___u2___expa[3'h7+:32'h00000001]) & fpu___u2___expb[3'h7+:32'h00000001]);
	assign fpu___u2___exp_ovf_d[1'h1+:32'h00000001] = (fpu___u2___op_div ? fpu___u2___co2 : ((~fpu___u2___expa[3'h7+:32'h00000001] & ~fpu___u2___expb[3'h7+:32'h00000001]) & fpu___u2___exp_tmp2[3'h7+:32'h00000001]) | fpu___u2___co2);
	always @(posedge clk) fpu___exp_ovf <= fpu___u2___exp_ovf_d;
	assign fpu___u2___underflow_d[2'h0+:32'h00000001] = ((8'h7f > fpu___u2___exp_tmp1) & ~fpu___u2___co1) & ~(((fpu___u2___opa_00 | fpu___u2___opb_00) | fpu___u2___expa_dn) | fpu___u2___expb_dn);
	assign fpu___u2___underflow_d[2'h1+:32'h00000001] = ((((fpu___u2___expa[3'h7+:32'h00000001] | fpu___u2___expb[3'h7+:32'h00000001]) & ~fpu___u2___opa_00) & ~fpu___u2___opb_00) | (fpu___u2___expa_dn & ~fpu___u2___fracta_00)) | (fpu___u2___expb_dn & ~fpu___u2___fractb_00);
	assign fpu___u2___underflow_d[2'h2+:32'h00000001] = (~fpu___u2___opa_00 & ~fpu___u2___opb_00) & (8'h7f == fpu___u2___exp_tmp1);
	always @(posedge clk) fpu___underflow_fmul_d <= fpu___u2___underflow_d;
	always @(posedge clk) fpu___inf_mul <= (fpu___u2___op_div ? fpu___u2___expb_dn & ~fpu___u2___expa[3'h7+:32'h00000001] : 9'h17e < {fpu___u2___co1, fpu___u2___exp_tmp1});
	always @(fpu___u2___signa or fpu___u2___signb)
		case ({fpu___u2___signa, fpu___u2___signb})
			2'h0: fpu___u2___sign_d = 1'h0;
			2'h1: fpu___u2___sign_d = 1'h1;
			2'h2: fpu___u2___sign_d = 1'h1;
			2'h3: fpu___u2___sign_d = 1'h0;
		endcase
	always @(posedge clk) fpu___sign_mul <= fpu___u2___sign_d;
	always @(posedge clk) fpu___sign_exe <= fpu___u2___signa & fpu___u2___signb;
	assign fpu___u3___add = fpu___fasu_op;
	assign fpu___u3___opa = fpu___fracta;
	assign fpu___u3___opb = fpu___fractb;
	assign fpu___u3___sum = fpu___fract_out_d;
	assign fpu___u3___co = fpu___co_d;
	assign ___sel_temp_9 = (fpu___fasu_op ? {1'b0, fpu___fracta} + {1'b0, fpu___fractb} : {1'b0, fpu___fracta} - {1'b0, fpu___fractb});
	assign fpu___co_d = ___sel_temp_9[32'h0000001b+:32'h00000001];
	assign ___sel_temp_10 = (fpu___fasu_op ? {1'b0, fpu___fracta} + {1'b0, fpu___fractb} : {1'b0, fpu___fracta} - {1'b0, fpu___fractb});
	assign fpu___fract_out_d = ___sel_temp_10[32'h00000000+:32'h0000001b];
	assign fpu___u5___clk = fpu___clk;
	assign fpu___u5___opa = fpu___fracta_mul;
	assign fpu___u5___opb = fpu___fractb_mul;
	wire [48:1] sv2v_tmp_6956B;
	assign sv2v_tmp_6956B = fpu___prod;
	always @(*) fpu___u5___prod = sv2v_tmp_6956B;
	always @(posedge clk) fpu___u5___prod1 <= {24'b000000000000000000000000, fpu___fracta_mul} * {24'b000000000000000000000000, fpu___fractb_mul};
	always @(posedge clk) fpu___prod <= fpu___u5___prod1;
	assign fpu___u_divider___clk = fpu___clk;
	assign fpu___u_divider___dividend = fpu___fdiv_opa;
	assign fpu___u_divider___divisor = fpu___fractb_mul;
	assign fpu___u_divider___merchant = fpu___quo;
	assign fpu___u_divider___remainder = fpu_____Vcellout__u_divider__remainder;
	assign fpu___u_divider___remainder_t1[5'h10] = fpu___u_divider_____Vcellout__u_divider_step0__remainder;
	assign fpu___u_divider___merchant_t1[5'h10] = fpu___u_divider_____Vcellout__u_divider_step0__merchant;
	assign fpu___u_divider___divisor_t1[5'h10] = fpu___u_divider_____Vcellout__u_divider_step0__divisor_kp;
	assign fpu___u_divider___dividend_t1[5'h10] = fpu___u_divider_____Vcellout__u_divider_step0__dividend_kp;
	assign fpu___u_divider_____Vcellinp__u_divider_step0__dividend_ci = fpu___fdiv_opa[6'h00+:32'h00000031];
	assign fpu___u_divider_____Vcellinp__u_divider_step0__dividend = {24'b000000000000000000000000, fpu___fdiv_opa[6'h31+:32'h00000001]};
	always @(posedge clk) begin
		fpu___u_divider___dividend_t2_r <= fpu___u_divider___dividend_t1[5'h00];
		fpu___u_divider___divisor_t2_r <= fpu___u_divider___divisor_t1[5'h00];
		fpu___u_divider___merchant_t2_r <= fpu___u_divider___merchant_t1[5'h00];
		fpu___u_divider___remainder_t2_r <= fpu___u_divider___remainder_t1[5'h00];
	end
	assign fpu___u_divider___dividend_t2[5'h10] = fpu___u_divider___dividend_t2_r;
	assign fpu___u_divider___divisor_t2[5'h10] = fpu___u_divider___divisor_t2_r;
	assign fpu___u_divider___merchant_t2[5'h10] = fpu___u_divider___merchant_t2_r;
	assign fpu___u_divider___remainder_t2[5'h10] = fpu___u_divider___remainder_t2_r;
	always @(posedge clk) begin
		fpu___u_divider___dividend_t3_r <= fpu___u_divider___dividend_t2[5'h00];
		fpu___u_divider___divisor_t3_r <= fpu___u_divider___divisor_t2[5'h00];
		fpu___u_divider___merchant_t3_r <= fpu___u_divider___merchant_t2[5'h00];
		fpu___u_divider___remainder_t3_r <= fpu___u_divider___remainder_t2[5'h00];
	end
	assign fpu___u_divider___dividend_t3[5'h11] = fpu___u_divider___dividend_t3_r;
	assign fpu___u_divider___divisor_t3[5'h11] = fpu___u_divider___divisor_t3_r;
	assign fpu___u_divider___merchant_t3[5'h11] = fpu___u_divider___merchant_t3_r;
	assign fpu___u_divider___remainder_t3[5'h11] = fpu___u_divider___remainder_t3_r;
	assign fpu___quo = fpu___u_divider___merchant_t3[5'h00];
	assign fpu_____Vcellout__u_divider__remainder = fpu___u_divider___remainder_t3[5'h00];
	assign fpu___u_divider___remainder_t1[5'h0f] = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h0f] = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h0f] = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h0f] = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h10], fpu___u_divider___dividend_t1[5'h10][6'h30+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h0e] = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h0e] = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h0e] = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h0e] = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h0f], fpu___u_divider___dividend_t1[5'h0f][6'h2f+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h0d] = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h0d] = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h0d] = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h0d] = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h0e], fpu___u_divider___dividend_t1[5'h0e][6'h2e+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h0c] = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h0c] = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h0c] = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h0c] = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h0d], fpu___u_divider___dividend_t1[5'h0d][6'h2d+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h0b] = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h0b] = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h0b] = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h0b] = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h0c], fpu___u_divider___dividend_t1[5'h0c][6'h2c+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h0a] = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h0a] = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h0a] = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h0a] = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h0b], fpu___u_divider___dividend_t1[5'h0b][6'h2b+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h09] = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h09] = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h09] = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h09] = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h0a], fpu___u_divider___dividend_t1[5'h0a][6'h2a+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h08] = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h08] = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h08] = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h08] = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h09], fpu___u_divider___dividend_t1[5'h09][6'h29+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h07] = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h07] = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h07] = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h07] = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h08], fpu___u_divider___dividend_t1[5'h08][6'h28+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h06] = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h06] = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h06] = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h06] = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h07], fpu___u_divider___dividend_t1[5'h07][6'h27+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h05] = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h05] = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h05] = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h05] = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h06], fpu___u_divider___dividend_t1[5'h06][6'h26+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h04] = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h04] = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h04] = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h04] = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h05], fpu___u_divider___dividend_t1[5'h05][6'h25+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h03] = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h03] = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h03] = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h03] = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h04], fpu___u_divider___dividend_t1[5'h04][6'h24+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h02] = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h02] = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h02] = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h02] = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h03], fpu___u_divider___dividend_t1[5'h03][6'h23+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h01] = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h01] = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h01] = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h01] = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h02], fpu___u_divider___dividend_t1[5'h02][6'h22+:32'h00000001]};
	assign fpu___u_divider___remainder_t1[5'h00] = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__remainder;
	assign fpu___u_divider___merchant_t1[5'h00] = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__merchant;
	assign fpu___u_divider___dividend_t1[5'h00] = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__dividend_kp;
	assign fpu___u_divider___divisor_t1[5'h00] = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend_ci = fpu___u_divider___dividend_t1[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__merchant_ci = fpu___u_divider___merchant_t1[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__divisor = fpu___u_divider___divisor_t1[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend = {fpu___u_divider___remainder_t1[5'h01], fpu___u_divider___dividend_t1[5'h01][6'h21+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h0f] = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h0f] = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h0f] = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h0f] = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h10], fpu___u_divider___dividend_t2[5'h10][6'h20+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h0e] = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h0e] = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h0e] = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h0e] = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h0f], fpu___u_divider___dividend_t2[5'h0f][6'h1f+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h0d] = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h0d] = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h0d] = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h0d] = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h0e], fpu___u_divider___dividend_t2[5'h0e][6'h1e+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h0c] = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h0c] = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h0c] = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h0c] = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h0d], fpu___u_divider___dividend_t2[5'h0d][6'h1d+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h0b] = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h0b] = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h0b] = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h0b] = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h0c], fpu___u_divider___dividend_t2[5'h0c][6'h1c+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h0a] = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h0a] = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h0a] = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h0a] = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h0b], fpu___u_divider___dividend_t2[5'h0b][6'h1b+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h09] = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h09] = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h09] = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h09] = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h0a], fpu___u_divider___dividend_t2[5'h0a][6'h1a+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h08] = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h08] = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h08] = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h08] = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h09], fpu___u_divider___dividend_t2[5'h09][6'h19+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h07] = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h07] = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h07] = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h07] = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h08], fpu___u_divider___dividend_t2[5'h08][6'h18+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h06] = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h06] = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h06] = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h06] = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h07], fpu___u_divider___dividend_t2[5'h07][6'h17+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h05] = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h05] = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h05] = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h05] = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h06], fpu___u_divider___dividend_t2[5'h06][6'h16+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h04] = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h04] = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h04] = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h04] = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h05], fpu___u_divider___dividend_t2[5'h05][6'h15+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h03] = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h03] = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h03] = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h03] = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h04], fpu___u_divider___dividend_t2[5'h04][6'h14+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h02] = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h02] = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h02] = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h02] = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h03], fpu___u_divider___dividend_t2[5'h03][6'h13+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h01] = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h01] = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h01] = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h01] = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h02], fpu___u_divider___dividend_t2[5'h02][6'h12+:32'h00000001]};
	assign fpu___u_divider___remainder_t2[5'h00] = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__remainder;
	assign fpu___u_divider___merchant_t2[5'h00] = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__merchant;
	assign fpu___u_divider___dividend_t2[5'h00] = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__dividend_kp;
	assign fpu___u_divider___divisor_t2[5'h00] = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend_ci = fpu___u_divider___dividend_t2[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__merchant_ci = fpu___u_divider___merchant_t2[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__divisor = fpu___u_divider___divisor_t2[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend = {fpu___u_divider___remainder_t2[5'h01], fpu___u_divider___dividend_t2[5'h01][6'h11+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h10] = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h10] = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h10] = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h10] = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h11];
	assign fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h11];
	assign fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h11];
	assign fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h11], fpu___u_divider___dividend_t3[5'h11][6'h10+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h0f] = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h0f] = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h0f] = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h0f] = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h10];
	assign fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h10], fpu___u_divider___dividend_t3[5'h10][6'h0f+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h0e] = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h0e] = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h0e] = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h0e] = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h0f];
	assign fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h0f], fpu___u_divider___dividend_t3[5'h0f][6'h0e+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h0d] = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h0d] = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h0d] = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h0d] = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h0e];
	assign fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h0e], fpu___u_divider___dividend_t3[5'h0e][6'h0d+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h0c] = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h0c] = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h0c] = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h0c] = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h0d];
	assign fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h0d], fpu___u_divider___dividend_t3[5'h0d][6'h0c+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h0b] = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h0b] = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h0b] = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h0b] = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h0c];
	assign fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h0c], fpu___u_divider___dividend_t3[5'h0c][6'h0b+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h0a] = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h0a] = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h0a] = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h0a] = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h0b];
	assign fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h0b], fpu___u_divider___dividend_t3[5'h0b][6'h0a+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h09] = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h09] = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h09] = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h09] = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h0a];
	assign fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h0a], fpu___u_divider___dividend_t3[5'h0a][6'h09+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h08] = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h08] = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h08] = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h08] = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h09];
	assign fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h09], fpu___u_divider___dividend_t3[5'h09][6'h08+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h07] = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h07] = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h07] = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h07] = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h08];
	assign fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h08], fpu___u_divider___dividend_t3[5'h08][6'h07+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h06] = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h06] = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h06] = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h06] = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h07];
	assign fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h07], fpu___u_divider___dividend_t3[5'h07][6'h06+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h05] = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h05] = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h05] = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h05] = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h06];
	assign fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h06], fpu___u_divider___dividend_t3[5'h06][6'h05+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h04] = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h04] = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h04] = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h04] = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h05];
	assign fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h05], fpu___u_divider___dividend_t3[5'h05][6'h04+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h03] = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h03] = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h03] = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h03] = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h04];
	assign fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h04], fpu___u_divider___dividend_t3[5'h04][6'h03+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h02] = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h02] = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h02] = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h02] = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h03];
	assign fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h03], fpu___u_divider___dividend_t3[5'h03][6'h02+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h01] = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h01] = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h01] = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h01] = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h02];
	assign fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h02], fpu___u_divider___dividend_t3[5'h02][6'h01+:32'h00000001]};
	assign fpu___u_divider___remainder_t3[5'h00] = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__remainder;
	assign fpu___u_divider___merchant_t3[5'h00] = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__merchant;
	assign fpu___u_divider___dividend_t3[5'h00] = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__dividend_kp;
	assign fpu___u_divider___divisor_t3[5'h00] = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__divisor_kp;
	assign fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend_ci = fpu___u_divider___dividend_t3[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__merchant_ci = fpu___u_divider___merchant_t3[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__divisor = fpu___u_divider___divisor_t3[5'h01];
	assign fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend = {fpu___u_divider___remainder_t3[5'h01], fpu___u_divider___dividend_t3[5'h01][6'h00+:32'h00000001]};
	assign fpu___u_divider___u_divider_step0___dividend = fpu___u_divider_____Vcellinp__u_divider_step0__dividend;
	assign fpu___u_divider___u_divider_step0___divisor = fpu___u_divider___divisor;
	assign fpu___u_divider___u_divider_step0___dividend_ci = fpu___u_divider_____Vcellinp__u_divider_step0__dividend_ci;
	assign fpu___u_divider___u_divider_step0___dividend_kp = fpu___u_divider_____Vcellout__u_divider_step0__dividend_kp;
	assign fpu___u_divider___u_divider_step0___divisor_kp = fpu___u_divider_____Vcellout__u_divider_step0__divisor_kp;
	assign fpu___u_divider___u_divider_step0___merchant = fpu___u_divider_____Vcellout__u_divider_step0__merchant;
	assign fpu___u_divider___u_divider_step0___remainder = fpu___u_divider_____Vcellout__u_divider_step0__remainder;
	assign fpu___u_divider_____Vcellout__u_divider_step0__divisor_kp = fpu___fractb_mul;
	assign fpu___u_divider_____Vcellout__u_divider_step0__dividend_kp = fpu___u_divider_____Vcellinp__u_divider_step0__dividend_ci;
	assign fpu___u_divider___u_divider_step0___geq = fpu___u_divider_____Vcellinp__u_divider_step0__dividend >= {1'b0, fpu___fractb_mul};
	assign fpu___u_divider_____Vcellout__u_divider_step0__merchant = (fpu___u_divider___u_divider_step0___geq ? 50'h0000000000001 : 50'h0000000000000);
	assign ___sel_temp_11 = (fpu___u_divider___u_divider_step0___geq ? fpu___u_divider_____Vcellinp__u_divider_step0__dividend - {1'b0, fpu___fractb_mul} : fpu___u_divider_____Vcellinp__u_divider_step0__dividend);
	assign fpu___u_divider_____Vcellout__u_divider_step0__remainder = ___sel_temp_11[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part11___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part11___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part11___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part11___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part11___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part11___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part11___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part11___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part11___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__merchant = (fpu___u_divider___gen_part11___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_12 = (fpu___u_divider___gen_part11___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part11___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part11___u_divider_step1__remainder = ___sel_temp_12[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part12___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part12___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part12___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part12___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part12___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part12___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part12___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part12___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part12___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__merchant = (fpu___u_divider___gen_part12___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_13 = (fpu___u_divider___gen_part12___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part12___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part12___u_divider_step1__remainder = ___sel_temp_13[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part13___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part13___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part13___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part13___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part13___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part13___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part13___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part13___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part13___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__merchant = (fpu___u_divider___gen_part13___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_14 = (fpu___u_divider___gen_part13___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part13___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part13___u_divider_step1__remainder = ___sel_temp_14[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part14___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part14___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part14___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part14___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part14___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part14___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part14___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part14___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part14___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__merchant = (fpu___u_divider___gen_part14___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_15 = (fpu___u_divider___gen_part14___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part14___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part14___u_divider_step1__remainder = ___sel_temp_15[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part15___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part15___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part15___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part15___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part15___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part15___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part15___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part15___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part15___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__merchant = (fpu___u_divider___gen_part15___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_16 = (fpu___u_divider___gen_part15___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part15___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part15___u_divider_step1__remainder = ___sel_temp_16[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part16___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part16___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part16___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part16___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part16___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part16___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part16___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part16___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part16___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__merchant = (fpu___u_divider___gen_part16___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_17 = (fpu___u_divider___gen_part16___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part16___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part16___u_divider_step1__remainder = ___sel_temp_17[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part17___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part17___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part17___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part17___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part17___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part17___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part17___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part17___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part17___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__merchant = (fpu___u_divider___gen_part17___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_18 = (fpu___u_divider___gen_part17___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part17___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part17___u_divider_step1__remainder = ___sel_temp_18[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part18___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part18___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part18___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part18___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part18___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part18___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part18___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part18___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part18___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__merchant = (fpu___u_divider___gen_part18___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_19 = (fpu___u_divider___gen_part18___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part18___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part18___u_divider_step1__remainder = ___sel_temp_19[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part19___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part19___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part19___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part19___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part19___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part19___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part19___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part19___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part19___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__merchant = (fpu___u_divider___gen_part19___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_20 = (fpu___u_divider___gen_part19___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part19___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part19___u_divider_step1__remainder = ___sel_temp_20[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part110___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part110___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part110___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part110___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part110___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part110___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part110___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part110___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part110___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__merchant = (fpu___u_divider___gen_part110___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_21 = (fpu___u_divider___gen_part110___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part110___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part110___u_divider_step1__remainder = ___sel_temp_21[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part111___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part111___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part111___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part111___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part111___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part111___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part111___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part111___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part111___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__merchant = (fpu___u_divider___gen_part111___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_22 = (fpu___u_divider___gen_part111___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part111___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part111___u_divider_step1__remainder = ___sel_temp_22[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part112___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part112___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part112___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part112___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part112___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part112___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part112___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part112___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part112___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__merchant = (fpu___u_divider___gen_part112___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_23 = (fpu___u_divider___gen_part112___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part112___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part112___u_divider_step1__remainder = ___sel_temp_23[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part113___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part113___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part113___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part113___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part113___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part113___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part113___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part113___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part113___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__merchant = (fpu___u_divider___gen_part113___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_24 = (fpu___u_divider___gen_part113___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part113___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part113___u_divider_step1__remainder = ___sel_temp_24[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part114___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part114___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part114___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part114___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part114___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part114___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part114___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part114___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part114___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__merchant = (fpu___u_divider___gen_part114___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_25 = (fpu___u_divider___gen_part114___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part114___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part114___u_divider_step1__remainder = ___sel_temp_25[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part115___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part115___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part115___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part115___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part115___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part115___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part115___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part115___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part115___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__merchant = (fpu___u_divider___gen_part115___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_26 = (fpu___u_divider___gen_part115___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part115___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part115___u_divider_step1__remainder = ___sel_temp_26[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part116___u_divider_step1___dividend = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend;
	assign fpu___u_divider___gen_part116___u_divider_step1___divisor = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__divisor;
	assign fpu___u_divider___gen_part116___u_divider_step1___merchant_ci = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__merchant_ci;
	assign fpu___u_divider___gen_part116___u_divider_step1___dividend_ci = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part116___u_divider_step1___dividend_kp = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__dividend_kp;
	assign fpu___u_divider___gen_part116___u_divider_step1___divisor_kp = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__divisor_kp;
	assign fpu___u_divider___gen_part116___u_divider_step1___merchant = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__merchant;
	assign fpu___u_divider___gen_part116___u_divider_step1___remainder = fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__remainder;
	assign fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__divisor_kp = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__divisor;
	assign fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__dividend_kp = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend_ci;
	assign fpu___u_divider___gen_part116___u_divider_step1___geq = fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__divisor};
	assign fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__merchant = (fpu___u_divider___gen_part116___u_divider_step1___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__merchant_ci << 32'sh00000001);
	assign ___sel_temp_27 = (fpu___u_divider___gen_part116___u_divider_step1___geq ? fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__divisor} : fpu___u_divider_____Vcellinp__gen_part116___u_divider_step1__dividend);
	assign fpu___u_divider_____Vcellout__gen_part116___u_divider_step1__remainder = ___sel_temp_27[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part21___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part21___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part21___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part21___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part21___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part21___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part21___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part21___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part21___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__merchant = (fpu___u_divider___gen_part21___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_28 = (fpu___u_divider___gen_part21___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part21___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part21___u_divider_step2__remainder = ___sel_temp_28[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part22___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part22___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part22___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part22___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part22___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part22___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part22___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part22___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part22___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__merchant = (fpu___u_divider___gen_part22___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_29 = (fpu___u_divider___gen_part22___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part22___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part22___u_divider_step2__remainder = ___sel_temp_29[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part23___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part23___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part23___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part23___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part23___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part23___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part23___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part23___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part23___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__merchant = (fpu___u_divider___gen_part23___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_30 = (fpu___u_divider___gen_part23___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part23___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part23___u_divider_step2__remainder = ___sel_temp_30[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part24___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part24___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part24___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part24___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part24___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part24___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part24___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part24___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part24___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__merchant = (fpu___u_divider___gen_part24___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_31 = (fpu___u_divider___gen_part24___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part24___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part24___u_divider_step2__remainder = ___sel_temp_31[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part25___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part25___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part25___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part25___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part25___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part25___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part25___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part25___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part25___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__merchant = (fpu___u_divider___gen_part25___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_32 = (fpu___u_divider___gen_part25___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part25___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part25___u_divider_step2__remainder = ___sel_temp_32[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part26___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part26___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part26___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part26___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part26___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part26___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part26___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part26___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part26___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__merchant = (fpu___u_divider___gen_part26___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_33 = (fpu___u_divider___gen_part26___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part26___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part26___u_divider_step2__remainder = ___sel_temp_33[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part27___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part27___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part27___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part27___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part27___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part27___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part27___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part27___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part27___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__merchant = (fpu___u_divider___gen_part27___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_34 = (fpu___u_divider___gen_part27___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part27___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part27___u_divider_step2__remainder = ___sel_temp_34[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part28___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part28___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part28___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part28___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part28___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part28___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part28___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part28___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part28___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__merchant = (fpu___u_divider___gen_part28___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_35 = (fpu___u_divider___gen_part28___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part28___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part28___u_divider_step2__remainder = ___sel_temp_35[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part29___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part29___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part29___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part29___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part29___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part29___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part29___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part29___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part29___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__merchant = (fpu___u_divider___gen_part29___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_36 = (fpu___u_divider___gen_part29___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part29___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part29___u_divider_step2__remainder = ___sel_temp_36[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part210___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part210___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part210___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part210___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part210___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part210___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part210___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part210___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part210___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__merchant = (fpu___u_divider___gen_part210___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_37 = (fpu___u_divider___gen_part210___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part210___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part210___u_divider_step2__remainder = ___sel_temp_37[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part211___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part211___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part211___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part211___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part211___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part211___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part211___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part211___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part211___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__merchant = (fpu___u_divider___gen_part211___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_38 = (fpu___u_divider___gen_part211___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part211___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part211___u_divider_step2__remainder = ___sel_temp_38[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part212___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part212___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part212___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part212___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part212___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part212___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part212___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part212___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part212___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__merchant = (fpu___u_divider___gen_part212___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_39 = (fpu___u_divider___gen_part212___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part212___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part212___u_divider_step2__remainder = ___sel_temp_39[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part213___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part213___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part213___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part213___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part213___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part213___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part213___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part213___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part213___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__merchant = (fpu___u_divider___gen_part213___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_40 = (fpu___u_divider___gen_part213___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part213___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part213___u_divider_step2__remainder = ___sel_temp_40[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part214___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part214___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part214___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part214___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part214___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part214___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part214___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part214___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part214___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__merchant = (fpu___u_divider___gen_part214___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_41 = (fpu___u_divider___gen_part214___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part214___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part214___u_divider_step2__remainder = ___sel_temp_41[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part215___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part215___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part215___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part215___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part215___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part215___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part215___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part215___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part215___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__merchant = (fpu___u_divider___gen_part215___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_42 = (fpu___u_divider___gen_part215___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part215___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part215___u_divider_step2__remainder = ___sel_temp_42[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part216___u_divider_step2___dividend = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend;
	assign fpu___u_divider___gen_part216___u_divider_step2___divisor = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__divisor;
	assign fpu___u_divider___gen_part216___u_divider_step2___merchant_ci = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__merchant_ci;
	assign fpu___u_divider___gen_part216___u_divider_step2___dividend_ci = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part216___u_divider_step2___dividend_kp = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__dividend_kp;
	assign fpu___u_divider___gen_part216___u_divider_step2___divisor_kp = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__divisor_kp;
	assign fpu___u_divider___gen_part216___u_divider_step2___merchant = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__merchant;
	assign fpu___u_divider___gen_part216___u_divider_step2___remainder = fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__remainder;
	assign fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__divisor_kp = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__divisor;
	assign fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__dividend_kp = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend_ci;
	assign fpu___u_divider___gen_part216___u_divider_step2___geq = fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__divisor};
	assign fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__merchant = (fpu___u_divider___gen_part216___u_divider_step2___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__merchant_ci << 32'sh00000001);
	assign ___sel_temp_43 = (fpu___u_divider___gen_part216___u_divider_step2___geq ? fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__divisor} : fpu___u_divider_____Vcellinp__gen_part216___u_divider_step2__dividend);
	assign fpu___u_divider_____Vcellout__gen_part216___u_divider_step2__remainder = ___sel_temp_43[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part31___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part31___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part31___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part31___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part31___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part31___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part31___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part31___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part31___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__merchant = (fpu___u_divider___gen_part31___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_44 = (fpu___u_divider___gen_part31___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part31___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part31___u_divider_step3__remainder = ___sel_temp_44[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part32___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part32___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part32___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part32___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part32___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part32___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part32___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part32___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part32___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__merchant = (fpu___u_divider___gen_part32___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_45 = (fpu___u_divider___gen_part32___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part32___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part32___u_divider_step3__remainder = ___sel_temp_45[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part33___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part33___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part33___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part33___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part33___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part33___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part33___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part33___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part33___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__merchant = (fpu___u_divider___gen_part33___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_46 = (fpu___u_divider___gen_part33___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part33___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part33___u_divider_step3__remainder = ___sel_temp_46[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part34___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part34___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part34___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part34___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part34___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part34___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part34___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part34___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part34___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__merchant = (fpu___u_divider___gen_part34___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_47 = (fpu___u_divider___gen_part34___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part34___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part34___u_divider_step3__remainder = ___sel_temp_47[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part35___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part35___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part35___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part35___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part35___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part35___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part35___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part35___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part35___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__merchant = (fpu___u_divider___gen_part35___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_48 = (fpu___u_divider___gen_part35___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part35___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part35___u_divider_step3__remainder = ___sel_temp_48[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part36___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part36___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part36___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part36___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part36___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part36___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part36___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part36___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part36___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__merchant = (fpu___u_divider___gen_part36___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_49 = (fpu___u_divider___gen_part36___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part36___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part36___u_divider_step3__remainder = ___sel_temp_49[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part37___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part37___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part37___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part37___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part37___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part37___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part37___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part37___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part37___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__merchant = (fpu___u_divider___gen_part37___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_50 = (fpu___u_divider___gen_part37___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part37___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part37___u_divider_step3__remainder = ___sel_temp_50[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part38___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part38___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part38___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part38___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part38___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part38___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part38___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part38___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part38___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__merchant = (fpu___u_divider___gen_part38___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_51 = (fpu___u_divider___gen_part38___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part38___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part38___u_divider_step3__remainder = ___sel_temp_51[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part39___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part39___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part39___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part39___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part39___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part39___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part39___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part39___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part39___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__merchant = (fpu___u_divider___gen_part39___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_52 = (fpu___u_divider___gen_part39___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part39___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part39___u_divider_step3__remainder = ___sel_temp_52[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part310___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part310___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part310___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part310___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part310___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part310___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part310___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part310___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part310___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__merchant = (fpu___u_divider___gen_part310___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_53 = (fpu___u_divider___gen_part310___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part310___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part310___u_divider_step3__remainder = ___sel_temp_53[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part311___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part311___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part311___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part311___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part311___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part311___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part311___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part311___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part311___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__merchant = (fpu___u_divider___gen_part311___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_54 = (fpu___u_divider___gen_part311___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part311___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part311___u_divider_step3__remainder = ___sel_temp_54[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part312___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part312___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part312___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part312___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part312___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part312___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part312___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part312___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part312___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__merchant = (fpu___u_divider___gen_part312___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_55 = (fpu___u_divider___gen_part312___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part312___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part312___u_divider_step3__remainder = ___sel_temp_55[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part313___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part313___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part313___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part313___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part313___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part313___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part313___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part313___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part313___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__merchant = (fpu___u_divider___gen_part313___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_56 = (fpu___u_divider___gen_part313___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part313___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part313___u_divider_step3__remainder = ___sel_temp_56[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part314___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part314___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part314___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part314___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part314___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part314___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part314___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part314___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part314___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__merchant = (fpu___u_divider___gen_part314___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_57 = (fpu___u_divider___gen_part314___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part314___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part314___u_divider_step3__remainder = ___sel_temp_57[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part315___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part315___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part315___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part315___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part315___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part315___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part315___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part315___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part315___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__merchant = (fpu___u_divider___gen_part315___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_58 = (fpu___u_divider___gen_part315___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part315___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part315___u_divider_step3__remainder = ___sel_temp_58[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part316___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part316___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part316___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part316___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part316___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part316___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part316___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part316___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part316___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__merchant = (fpu___u_divider___gen_part316___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_59 = (fpu___u_divider___gen_part316___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part316___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part316___u_divider_step3__remainder = ___sel_temp_59[32'h00000000+:32'h00000018];
	assign fpu___u_divider___gen_part317___u_divider_step3___dividend = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend;
	assign fpu___u_divider___gen_part317___u_divider_step3___divisor = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__divisor;
	assign fpu___u_divider___gen_part317___u_divider_step3___merchant_ci = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__merchant_ci;
	assign fpu___u_divider___gen_part317___u_divider_step3___dividend_ci = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part317___u_divider_step3___dividend_kp = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__dividend_kp;
	assign fpu___u_divider___gen_part317___u_divider_step3___divisor_kp = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__divisor_kp;
	assign fpu___u_divider___gen_part317___u_divider_step3___merchant = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__merchant;
	assign fpu___u_divider___gen_part317___u_divider_step3___remainder = fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__remainder;
	assign fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__divisor_kp = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__divisor;
	assign fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__dividend_kp = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend_ci;
	assign fpu___u_divider___gen_part317___u_divider_step3___geq = fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend >= {1'b0, fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__divisor};
	assign fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__merchant = (fpu___u_divider___gen_part317___u_divider_step3___geq ? 50'h0000000000001 | (fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__merchant_ci << 32'sh00000001) : fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__merchant_ci << 32'sh00000001);
	assign ___sel_temp_60 = (fpu___u_divider___gen_part317___u_divider_step3___geq ? fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend - {1'b0, fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__divisor} : fpu___u_divider_____Vcellinp__gen_part317___u_divider_step3__dividend);
	assign fpu___u_divider_____Vcellout__gen_part317___u_divider_step3__remainder = ___sel_temp_60[32'h00000000+:32'h00000018];
	assign fpu___u4___clk = fpu___clk;
	assign fpu___u4___fpu_op = fpu___fpu_op_r3;
	assign fpu___u4___opas = fpu___opas_r2;
	assign fpu___u4___sign = fpu___sign;
	assign fpu___u4___rmode = fpu___rmode_r3;
	assign fpu___u4___fract_in = fpu___fract_denorm;
	assign fpu___u4___exp_in = fpu___exp_r;
	assign fpu___u4___exp_ovf = fpu___exp_ovf_r;
	assign fpu___u4___opa_dn = fpu___opa_dn;
	assign fpu___u4___opb_dn = fpu___opb_dn;
	assign fpu___u4___rem_00 = fpu___remainder_00;
	assign fpu___u4___div_opa_ldz = fpu___div_opa_ldz_r2;
	assign fpu___u4___output_zero = fpu_____Vcellinp__u4__output_zero;
	assign fpu___u4___out = fpu___out_d;
	assign fpu___u4___ine = fpu___ine_d;
	assign fpu___u4___overflow = fpu___overflow_d;
	assign fpu___u4___underflow = fpu___underflow_d;
	assign fpu___u4___f2i_out_sign = fpu___f2i_out_sign;
	assign fpu___u4___op_dn = fpu___opa_dn | fpu___opb_dn;
	assign fpu___u4___op_mul = 3'h2 == fpu___fpu_op_r3;
	assign fpu___u4___op_div = 3'h3 == fpu___fpu_op_r3;
	assign fpu___u4___op_i2f = 3'h4 == fpu___fpu_op_r3;
	assign fpu___u4___op_f2i = 3'h5 == fpu___fpu_op_r3;
	always @(fpu___fract_denorm)
		case (fpu___fract_denorm)
			48'b1zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h01;
			48'b01zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h02;
			48'b001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h03;
			48'b0001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h04;
			48'b00001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h05;
			48'b000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h06;
			48'b0000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h07;
			48'b00000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h08;
			48'b000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h09;
			48'b0000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h0a;
			48'b00000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h0b;
			48'b000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h0c;
			48'b0000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h0d;
			48'b00000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h0e;
			48'b000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h0f;
			48'b0000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h10;
			48'b00000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h11;
			48'b000000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h12;
			48'b0000000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h13;
			48'b00000000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h14;
			48'b000000000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h15;
			48'b0000000000000000000001zzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h16;
			48'b00000000000000000000001zzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h17;
			48'b000000000000000000000001zzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h18;
			48'b0000000000000000000000001zzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h19;
			48'b00000000000000000000000001zzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h1a;
			48'b000000000000000000000000001zzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h1b;
			48'b0000000000000000000000000001zzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h1c;
			48'b00000000000000000000000000001zzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h1d;
			48'b000000000000000000000000000001zzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h1e;
			48'b0000000000000000000000000000001zzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h1f;
			48'b00000000000000000000000000000001zzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h20;
			48'b000000000000000000000000000000001zzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h21;
			48'b0000000000000000000000000000000001zzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h22;
			48'b00000000000000000000000000000000001zzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h23;
			48'b000000000000000000000000000000000001zzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h24;
			48'b0000000000000000000000000000000000001zzzzzzzzzzz: fpu___u4___fi_ldz = 6'h25;
			48'b00000000000000000000000000000000000001zzzzzzzzzz: fpu___u4___fi_ldz = 6'h26;
			48'b000000000000000000000000000000000000001zzzzzzzzz: fpu___u4___fi_ldz = 6'h27;
			48'b0000000000000000000000000000000000000001zzzzzzzz: fpu___u4___fi_ldz = 6'h28;
			48'b00000000000000000000000000000000000000001zzzzzzz: fpu___u4___fi_ldz = 6'h29;
			48'b000000000000000000000000000000000000000001zzzzzz: fpu___u4___fi_ldz = 6'h2a;
			48'b0000000000000000000000000000000000000000001zzzzz: fpu___u4___fi_ldz = 6'h2b;
			48'b00000000000000000000000000000000000000000001zzzz: fpu___u4___fi_ldz = 6'h2c;
			48'b000000000000000000000000000000000000000000001zzz: fpu___u4___fi_ldz = 6'h2d;
			48'b0000000000000000000000000000000000000000000001zz: fpu___u4___fi_ldz = 6'h2e;
			48'b00000000000000000000000000000000000000000000001z: fpu___u4___fi_ldz = 6'h2f;
			48'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz: fpu___u4___fi_ldz = 6'h30;
		endcase
	assign fpu___u4___exp_in_ff = &fpu___exp_r;
	assign fpu___u4___exp_in_00 = ~(|fpu___exp_r);
	assign fpu___u4___exp_in_80 = fpu___exp_r[3'h7+:32'h00000001] & ~(|fpu___exp_r[3'h0+:32'h00000007]);
	assign fpu___u4___exp_out_ff = &fpu___u4___exp_out;
	assign fpu___u4___exp_out_00 = ~(|fpu___u4___exp_out);
	assign fpu___u4___exp_out_fe = &fpu___u4___exp_out[3'h1+:32'h00000007] & ~fpu___u4___exp_out[3'h0+:32'h00000001];
	assign fpu___u4___exp_out_final_ff = &fpu___u4___exp_out_final;
	assign fpu___u4___fract_out_7fffff = &fpu___u4___fract_out;
	assign fpu___u4___fract_out_00 = ~(|fpu___u4___fract_out);
	assign fpu___u4___fract_in_00 = ~(|fpu___fract_denorm);
	assign fpu___u4___rmode_00 = 2'h0 == fpu___rmode_r3;
	assign fpu___u4___rmode_01 = 2'h1 == fpu___rmode_r3;
	assign fpu___u4___rmode_10 = 2'h2 == fpu___rmode_r3;
	assign fpu___u4___rmode_11 = 2'h3 == fpu___rmode_r3;
	assign fpu___u4___dn = (~fpu___u4___op_mul & ~fpu___u4___op_div) & (fpu___u4___exp_in_00 | (fpu___u4___exp_next_mi[4'h8+:32'h00000001] & ~fpu___fract_denorm[6'h2f+:32'h00000001]));
	assign fpu___u4___fract_out_pl1 = 24'h000001 + {9'b000000000, fpu___u4___fract_out}[32'h00000000+:32'h00000018];
	assign fpu___u4___f2i_emin = (fpu___u4___rmode_00 ? 8'h7e : 8'h7f);
	assign fpu___u4___f2i_zero = ((~fpu___opas_r2 & (fpu___exp_r < fpu___u4___f2i_emin)) | (fpu___opas_r2 & (8'h9d < fpu___exp_r))) | ((fpu___opas_r2 & (fpu___exp_r < fpu___u4___f2i_emin)) & (fpu___u4___fract_in_00 | ~fpu___u4___rmode_11));
	assign fpu___u4___f2i_max = (~fpu___opas_r2 & (8'h9d < fpu___exp_r)) | (((fpu___opas_r2 & (fpu___exp_r < fpu___u4___f2i_emin)) & ~fpu___u4___fract_in_00) & fpu___u4___rmode_11);
	assign ___sel_temp_61 = (~fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___u4___exp_in_00 ? {1'b0, fpu___u4___exp_out} : fpu___u4___exp_in_mi1);
	assign fpu___u4___shft_co = ___sel_temp_61[32'h00000008+:32'h00000001];
	assign ___sel_temp_62 = (~fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___u4___exp_in_00 ? {1'b0, fpu___u4___exp_out} : fpu___u4___exp_in_mi1);
	assign fpu___u4___shftr_mul = ___sel_temp_62[32'h00000000+:32'h00000008];
	assign ___sel_temp_63 = (fpu___u4___exp_in_00 ? {4'b0000, fpu___div_opa_ldz_r2} : fpu___u4___div_scht1a);
	assign fpu___u4___div_shft1_co = ___sel_temp_63[32'h00000008+:32'h00000001];
	assign ___sel_temp_64 = (fpu___u4___exp_in_00 ? {4'b0000, fpu___div_opa_ldz_r2} : fpu___u4___div_scht1a);
	assign fpu___u4___div_shft1 = ___sel_temp_64[32'h00000000+:32'h00000008];
	assign fpu___u4___div_scht1a = {1'b0, fpu___exp_r} - {4'b0000, fpu___div_opa_ldz_r2};
	assign fpu___u4___div_shft2 = 8'h02 + fpu___exp_r;
	assign fpu___u4___div_shft3 = {3'b000, fpu___div_opa_ldz_r2} + fpu___exp_r;
	assign fpu___u4___div_shft4 = {3'b000, fpu___div_opa_ldz_r2} - fpu___exp_r;
	assign fpu___u4___div_dn = fpu___u4___op_dn & fpu___u4___div_shft1_co;
	assign fpu___u4___div_nr = ((fpu___u4___op_dn & fpu___exp_ovf_r[1'h1+:32'h00000001]) & ~(|fpu___fract_denorm[6'h17+:32'h00000018])) & (8'h16 < fpu___u4___div_shft3);
	assign fpu___u4___f2i_shft = fpu___exp_r - 8'h7d;
	assign ___sel_temp_65 = (fpu___u4___op_div ? {31'b0000000000000000000000000000000, fpu___u4___lr_div} : (fpu___u4___op_mul ? {31'b0000000000000000000000000000000, fpu___u4___lr_mul} : 32'sh00000001));
	assign fpu___u4___left_right = ___sel_temp_65[32'h00000000+:32'h00000001];
	assign ___sel_temp_66 = ((fpu___u4___op_dn & ~fpu___exp_ovf_r[1'h1+:32'h00000001]) & fpu___exp_ovf_r[1'h0+:32'h00000001] ? 32'sh00000001 : (fpu___u4___op_dn & fpu___exp_ovf_r[1'h1+:32'h00000001] ? 32'sh00000000 : (fpu___u4___op_dn & fpu___u4___div_shft1_co ? 32'sh00000000 : (fpu___u4___op_dn & fpu___u4___exp_out_00 ? 32'sh00000001 : ((~fpu___u4___op_dn & fpu___u4___exp_out_00) & ~fpu___exp_ovf_r[1'h1+:32'h00000001] ? 32'sh00000001 : (fpu___exp_ovf_r[1'h1+:32'h00000001] ? 32'sh00000000 : 32'sh00000001))))));
	assign fpu___u4___lr_div = ___sel_temp_66[32'h00000000+:32'h00000001];
	assign ___sel_temp_67 = ((fpu___u4___shft_co | (~fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___u4___exp_in_00)) | ((~fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___u4___exp_in_00) & (fpu___u4___exp_out1_co | fpu___u4___exp_out_00)) ? 32'sh00000001 : (fpu___exp_ovf_r[1'h1+:32'h00000001] | fpu___u4___exp_in_00 ? 32'sh00000000 : 32'sh00000001));
	assign fpu___u4___lr_mul = ___sel_temp_67[32'h00000000+:32'h00000001];
	assign fpu___u4___fasu_shift = (fpu___u4___dn | fpu___u4___exp_out_00 ? (fpu___u4___exp_in_00 ? 8'h02 : fpu___u4___exp_in_pl1[4'h0+:32'h00000008]) : {2'b00, fpu___u4___fi_ldz});
	assign fpu___u4___shift_right = (fpu___u4___op_div ? fpu___u4___shftr_div : fpu___u4___shftr_mul);
	assign fpu___u4___conv_shft = (fpu___u4___op_f2i ? fpu___u4___f2i_shft : {2'b00, fpu___u4___fi_ldz});
	assign fpu___u4___shift_left = (fpu___u4___op_div ? fpu___u4___shftl_div : (fpu___u4___op_mul ? fpu___u4___shftl_mul : (fpu___u4___op_f2i | fpu___u4___op_i2f ? fpu___u4___conv_shft : fpu___u4___fasu_shift)));
	assign fpu___u4___shftl_mul = ((fpu___u4___shft_co | (~fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___u4___exp_in_00)) | ((~fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___u4___exp_in_00) & (fpu___u4___exp_out1_co | fpu___u4___exp_out_00)) ? fpu___u4___exp_in_pl1[4'h0+:32'h00000008] : {2'b00, fpu___u4___fi_ldz});
	assign fpu___u4___shftl_div = ((fpu___u4___op_dn & fpu___u4___exp_out_00) & ~(~fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___exp_ovf_r[1'h0+:32'h00000001]) ? fpu___u4___div_shft1 : ((~fpu___u4___op_dn & fpu___u4___exp_out_00) & ~fpu___exp_ovf_r[1'h1+:32'h00000001] ? fpu___exp_r : {2'b00, fpu___u4___fi_ldz}));
	assign fpu___u4___shftr_div = (fpu___u4___op_dn & fpu___exp_ovf_r[1'h1+:32'h00000001] ? fpu___u4___div_shft3 : (fpu___u4___op_dn & fpu___u4___div_shft1_co ? fpu___u4___div_shft4 : fpu___u4___div_shft2));
	assign fpu___u4___fract_in_shftr = (|fpu___u4___shift_right[3'h6+:32'h00000002] ? 48'h000000000000 : fpu___fract_denorm >> fpu___u4___shift_right[3'h0+:32'h00000006]);
	assign fpu___u4___fract_in_shftl = (|fpu___u4___shift_left[3'h6+:32'h00000002] | (fpu___u4___f2i_zero & fpu___u4___op_f2i) ? 48'h000000000000 : fpu___fract_denorm << fpu___u4___shift_left[3'h0+:32'h00000006]);
	assign ___sel_temp_68 = (fpu___u4___left_right ? fpu___u4___fract_in_shftl : fpu___u4___fract_in_shftr);
	assign fpu___u4___fract_out = ___sel_temp_68[32'h00000019+:32'h00000017];
	assign ___sel_temp_69 = (fpu___u4___left_right ? fpu___u4___fract_in_shftl : fpu___u4___fract_in_shftr);
	assign fpu___u4___fract_trunc = ___sel_temp_69[32'h00000000+:32'h00000019];
	assign fpu___u4___fi_ldz_mi1 = fpu___u4___fi_ldz - 6'h01;
	assign fpu___u4___fi_ldz_mi22 = fpu___u4___fi_ldz - 6'h16;
	assign fpu___u4___exp_out_pl1 = 8'h01 + fpu___u4___exp_out;
	assign fpu___u4___exp_out_mi1 = fpu___u4___exp_out - 8'h01;
	assign fpu___u4___exp_in_pl1 = 9'h001 + {24'b000000000000000000000000, fpu___exp_r}[32'h00000000+:32'h00000009];
	assign fpu___u4___exp_in_mi1 = {24'b000000000000000000000000, fpu___exp_r}[32'h00000000+:32'h00000009] - 9'h001;
	assign fpu___u4___exp_out1_mi1 = fpu___u4___exp_out1 - 8'h01;
	assign fpu___u4___exp_next_mi = fpu___u4___exp_in_pl1 - {3'b000, fpu___u4___fi_ldz_mi1};
	assign fpu___u4___exp_fix_diva = fpu___exp_r - {2'b00, fpu___u4___fi_ldz_mi22};
	assign fpu___u4___exp_fix_divb = fpu___exp_r - {2'b00, fpu___u4___fi_ldz_mi1};
	assign fpu___u4___exp_zero = (((fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) & fpu___u4___op_mul) & (~fpu___u4___exp_rnd_adj2a | ~fpu___rmode_r3[1'h1+:32'h00000001])) | (fpu___u4___op_mul & fpu___u4___exp_out1_co);
	assign ___sel_temp_70 = (fpu___fract_denorm[6'h2f+:32'h00000001] ? fpu___u4___exp_in_pl1 : fpu___u4___exp_next_mi);
	assign fpu___u4___exp_out1_co = ___sel_temp_70[32'h00000008+:32'h00000001];
	assign ___sel_temp_71 = (fpu___fract_denorm[6'h2f+:32'h00000001] ? fpu___u4___exp_in_pl1 : fpu___u4___exp_next_mi);
	assign fpu___u4___exp_out1 = ___sel_temp_71[32'h00000000+:32'h00000008];
	assign ___sel_temp_72 = (fpu___opas_r2 ? (fpu___exp_r < fpu___u4___f2i_emin ? 32'sh00000000 : (8'h9d < fpu___exp_r ? 32'sh00000001 : {31'b0000000000000000000000000000000, fpu___opas_r2})) : (fpu___exp_r < fpu___u4___f2i_emin ? 32'sh00000000 : (8'h9d < fpu___exp_r ? 32'sh00000000 : {31'b0000000000000000000000000000000, fpu___opas_r2})));
	assign fpu___f2i_out_sign = ___sel_temp_72[32'h00000000+:32'h00000001];
	assign ___sel_temp_73 = (fpu___u4___fract_in_00 ? (fpu___opas_r2 ? 32'h0000009e : 32'sh00000000) : 32'h0000009e - {26'b00000000000000000000000000, fpu___u4___fi_ldz});
	assign fpu___u4___exp_i2f = ___sel_temp_73[32'h00000000+:32'h00000008];
	assign fpu___u4___exp_f2i_1 = {{32'sh00000008 {fpu___fract_denorm[6'h2f+:32'h00000001]}}, fpu___fract_denorm} << fpu___u4___f2i_shft;
	assign ___sel_temp_74 = (fpu___u4___f2i_zero ? 32'sh00000000 : (fpu___u4___f2i_max ? 32'h000000ff : {24'b000000000000000000000000, fpu___u4___exp_f2i_1[6'h30+:32'h00000008]}));
	assign fpu___u4___exp_f2i = ___sel_temp_74[32'h00000000+:32'h00000008];
	assign fpu___u4___conv_exp = (fpu___u4___op_f2i ? fpu___u4___exp_f2i : fpu___u4___exp_i2f);
	assign fpu___u4___exp_out = (fpu___u4___op_div ? fpu___u4___exp_div : (fpu___u4___op_f2i | fpu___u4___op_i2f ? fpu___u4___conv_exp : (fpu___u4___exp_zero ? 8'h00 : (fpu___u4___dn ? {6'b000000, fpu___fract_denorm[6'h2e+:32'h00000002]} : fpu___u4___exp_out1))));
	assign fpu___u4___ldz_all = {2'b00, fpu___div_opa_ldz_r2} + {1'b0, fpu___u4___fi_ldz};
	assign fpu___u4___ldz_dif = fpu___u4___fi_ldz_2 - {3'b000, fpu___div_opa_ldz_r2};
	assign fpu___u4___fi_ldz_2a = 7'h17 - {1'b0, fpu___u4___fi_ldz};
	assign fpu___u4___fi_ldz_2 = {fpu___u4___fi_ldz_2a[3'h6+:32'h00000001], fpu___u4___fi_ldz_2a};
	assign fpu___u4___div_exp1 = fpu___u4___exp_in_mi1 + {1'b0, fpu___u4___fi_ldz_2};
	assign fpu___u4___div_exp2 = fpu___u4___exp_in_pl1[32'h00000000+:32'h00000008] - {2'b00, fpu___u4___ldz_all}[32'h00000000+:32'h00000008];
	assign fpu___u4___div_exp3 = fpu___exp_r + fpu___u4___ldz_dif;
	assign ___sel_temp_75 = (fpu___opa_dn & fpu___opb_dn ? {24'b000000000000000000000000, fpu___u4___div_exp3} : (fpu___opb_dn ? {24'b000000000000000000000000, fpu___u4___div_exp1[4'h0+:32'h00000008]} : (fpu___opa_dn & ~((fpu___exp_r < {3'b000, fpu___div_opa_ldz_r2}) | (8'hfe < fpu___u4___div_exp2)) ? {24'b000000000000000000000000, fpu___u4___div_exp2} : (fpu___opa_dn | (fpu___u4___exp_in_00 & ~fpu___exp_ovf_r[1'h1+:32'h00000001]) ? 32'sh00000000 : {24'b000000000000000000000000, fpu___u4___exp_out1_mi1}))));
	assign fpu___u4___exp_div = ___sel_temp_75[32'h00000000+:32'h00000008];
	assign fpu___u4___div_inf = (fpu___opb_dn & ~fpu___opa_dn) & (8'h7f > fpu___u4___div_exp1[4'h0+:32'h00000008]);
	assign fpu___u4___grs_sel_div = fpu___u4___op_div & (((fpu___exp_ovf_r[1'h1+:32'h00000001] | fpu___u4___div_dn) | fpu___u4___exp_out1_co) | fpu___u4___exp_out_00);
	assign fpu___u4___g = (fpu___u4___grs_sel_div ? fpu___u4___fract_out[5'h00+:32'h00000001] : fpu___u4___fract_out[5'h00+:32'h00000001]);
	assign fpu___u4___r = (fpu___u4___grs_sel_div ? fpu___u4___fract_trunc[5'h18+:32'h00000001] & ~fpu___u4___div_nr : fpu___u4___fract_trunc[5'h18+:32'h00000001]);
	assign fpu___u4___s = (fpu___u4___grs_sel_div ? |fpu___u4___fract_trunc : |fpu___u4___fract_trunc[5'h00+:32'h00000018] | (fpu___u4___fract_trunc[5'h18+:32'h00000001] & fpu___u4___op_div));
	assign fpu___u4___round = (fpu___u4___g & fpu___u4___r) | (fpu___u4___r & fpu___u4___s);
	assign ___sel_temp_76 = (fpu___u4___round ? fpu___u4___fract_out_pl1 : {1'b0, fpu___u4___fract_out});
	assign fpu___u4___exp_rnd_adj0 = ___sel_temp_76[32'h00000017+:32'h00000001];
	assign ___sel_temp_77 = (fpu___u4___round ? fpu___u4___fract_out_pl1 : {1'b0, fpu___u4___fract_out});
	assign fpu___u4___fract_out_rnd0 = ___sel_temp_77[32'h00000000+:32'h00000017];
	assign fpu___u4___exp_out_rnd0 = (fpu___u4___exp_rnd_adj0 ? fpu___u4___exp_out_pl1 : fpu___u4___exp_out);
	assign fpu___u4___ovf0 = (fpu___u4___exp_out_final_ff & ~fpu___u4___rmode_01) & ~fpu___u4___op_f2i;
	assign fpu___u4___fract_out_rnd1 = (((fpu___u4___exp_out_ff & ~fpu___u4___op_div) & ~fpu___u4___dn) & ~fpu___u4___op_f2i ? 23'h7fffff : fpu___u4___fract_out);
	assign fpu___u4___exp_fix_div = (6'h16 < fpu___u4___fi_ldz ? fpu___u4___exp_fix_diva : fpu___u4___exp_fix_divb);
	assign fpu___u4___exp_out_rnd1 = (((fpu___u4___g & fpu___u4___r) & fpu___u4___s) & fpu___u4___exp_in_ff ? (fpu___u4___op_div ? fpu___u4___exp_fix_div : fpu___u4___exp_next_mi[4'h0+:32'h00000008]) : (fpu___u4___exp_out_ff & ~fpu___u4___op_f2i ? fpu___exp_r : fpu___u4___exp_out));
	assign fpu___u4___ovf1 = fpu___u4___exp_out_ff & ~fpu___u4___dn;
	assign fpu___u4___r_sign = fpu___sign;
	assign fpu___u4___round2a = (~fpu___u4___exp_out_fe | ~fpu___u4___fract_out_7fffff) | (fpu___u4___exp_out_fe & fpu___u4___fract_out_7fffff);
	assign fpu___u4___round2_fasu = ((fpu___u4___r | fpu___u4___s) & ~fpu___u4___r_sign) & (~fpu___u4___exp_out[3'h7+:32'h00000001] | (fpu___u4___exp_out[3'h7+:32'h00000001] & fpu___u4___round2a));
	assign fpu___u4___round2_fmul = ~fpu___u4___r_sign & (((fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___u4___fract_in_00) & ((((~fpu___u4___exp_out1_co | fpu___u4___op_dn) & ((fpu___u4___r | fpu___u4___s) | (~fpu___remainder_00 & fpu___u4___op_div))) | fpu___u4___fract_out_00) | (~fpu___u4___op_dn & ~fpu___u4___op_div))) | (((fpu___u4___r | fpu___u4___s) | (~fpu___remainder_00 & fpu___u4___op_div)) & (((~fpu___exp_ovf_r[1'h1+:32'h00000001] & (fpu___u4___exp_in_80 | ~fpu___exp_ovf_r[1'h0+:32'h00000001])) | fpu___u4___op_div) | ((fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) & fpu___u4___exp_out1_co))));
	assign fpu___u4___round2_f2i = fpu___u4___rmode_10 & (((|fpu___fract_denorm[6'h00+:32'h00000018] & ~fpu___opas_r2) & (8'h80 > fpu___exp_r)) | (|fpu___u4___fract_trunc));
	assign fpu___u4___round2 = (fpu___u4___op_mul | fpu___u4___op_div ? fpu___u4___round2_fmul : (fpu___u4___op_f2i ? fpu___u4___round2_f2i : fpu___u4___round2_fasu));
	assign ___sel_temp_78 = (fpu___u4___round2 ? fpu___u4___fract_out_pl1 : {1'b0, fpu___u4___fract_out});
	assign fpu___u4___exp_rnd_adj2a = ___sel_temp_78[32'h00000017+:32'h00000001];
	assign ___sel_temp_79 = (fpu___u4___round2 ? fpu___u4___fract_out_pl1 : {1'b0, fpu___u4___fract_out});
	assign fpu___u4___fract_out_rnd2a = ___sel_temp_79[32'h00000000+:32'h00000017];
	assign fpu___u4___exp_out_rnd2a = (fpu___u4___exp_rnd_adj2a ? (fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___u4___op_mul ? fpu___u4___exp_out_mi1 : fpu___u4___exp_out_pl1) : fpu___u4___exp_out);
	assign fpu___u4___fract_out_rnd2 = ((((fpu___u4___r_sign & fpu___u4___exp_out_ff) & ~fpu___u4___op_div) & ~fpu___u4___dn) & ~fpu___u4___op_f2i ? 23'h7fffff : fpu___u4___fract_out_rnd2a);
	assign fpu___u4___exp_out_rnd2 = ((fpu___u4___r_sign & fpu___u4___exp_out_ff) & ~fpu___u4___op_f2i ? 8'hfe : fpu___u4___exp_out_rnd2a);
	always @(fpu___rmode_r3 or fpu___u4___exp_out_rnd0 or fpu___u4___exp_out_rnd1 or fpu___u4___exp_out_rnd2)
		case ({30'b000000000000000000000000000000, fpu___rmode_r3})
			32'sh00000000: fpu___u4___exp_out_rnd = fpu___u4___exp_out_rnd0;
			32'sh00000001: fpu___u4___exp_out_rnd = fpu___u4___exp_out_rnd1;
			32'sh00000002, 32'sh00000003: fpu___u4___exp_out_rnd = fpu___u4___exp_out_rnd2;
		endcase
	always @(fpu___rmode_r3 or fpu___u4___fract_out_rnd0 or fpu___u4___fract_out_rnd1 or fpu___u4___fract_out_rnd2)
		case ({30'b000000000000000000000000000000, fpu___rmode_r3})
			32'sh00000000: fpu___u4___fract_out_rnd = fpu___u4___fract_out_rnd0;
			32'sh00000001: fpu___u4___fract_out_rnd = fpu___u4___fract_out_rnd1;
			32'sh00000002, 32'sh00000003: fpu___u4___fract_out_rnd = fpu___u4___fract_out_rnd2;
		endcase
	assign fpu___u4___max_num = ((~fpu___u4___rmode_00 & (fpu___u4___op_mul | fpu___u4___op_div)) & ((fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___exp_ovf_r[1'h0+:32'h00000001]) | ((((~fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) & fpu___u4___exp_in_ff) & (8'h18 > fpu___u4___fi_ldz_2)) & (8'hfe != fpu___u4___exp_out)))) | (fpu___u4___op_div & ((fpu___u4___rmode_01 & ((fpu___u4___div_inf | (fpu___u4___exp_out_ff & ~fpu___exp_ovf_r[1'h1+:32'h00000001])) | (fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___exp_ovf_r[1'h0+:32'h00000001]))) | ((fpu___rmode_r3[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h1+:32'h00000001]) & (((((fpu___exp_ovf_r[1'h0+:32'h00000001] & fpu___u4___exp_in_ff) & fpu___u4___r_sign) & fpu___fract_denorm[6'h2f+:32'h00000001]) | (fpu___u4___r_sign & (((fpu___fract_denorm[6'h2f+:32'h00000001] & fpu___u4___div_inf) | (((fpu___exp_r[3'h7+:32'h00000001] & ~fpu___u4___exp_out_rnd[3'h7+:32'h00000001]) & ~fpu___u4___exp_in_80) & (8'h7f != fpu___u4___exp_out))) | (((((fpu___exp_r[3'h7+:32'h00000001] & fpu___u4___exp_out_rnd[3'h7+:32'h00000001]) & fpu___u4___r_sign) & fpu___u4___exp_out_ff) & fpu___u4___op_dn) & (9'h0fe < fpu___u4___div_exp1))))) | ((fpu___u4___exp_in_00 & fpu___u4___r_sign) & (fpu___u4___div_inf | ((fpu___u4___r_sign & fpu___u4___exp_out_ff) & (8'h18 > fpu___u4___fi_ldz_2))))))));
	assign fpu___u4___inf_out = ((((fpu___rmode_r3[1'h1+:32'h00000001] & (fpu___u4___op_mul | fpu___u4___op_div)) & ~fpu___u4___r_sign) & ((fpu___u4___exp_in_ff & ~fpu___u4___op_div) | ((fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___exp_ovf_r[1'h0+:32'h00000001]) & (fpu___u4___exp_in_00 | fpu___exp_r[3'h7+:32'h00000001])))) | ((fpu___u4___div_inf & fpu___u4___op_div) & ((fpu___u4___rmode_00 | ((((fpu___rmode_r3[1'h1+:32'h00000001] & ~fpu___u4___exp_in_ff) & ~fpu___exp_ovf_r[1'h1+:32'h00000001]) & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) & ~fpu___u4___r_sign)) | ((((fpu___rmode_r3[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h1+:32'h00000001]) & fpu___exp_ovf_r[1'h0+:32'h00000001]) & fpu___u4___exp_in_00) & ~fpu___u4___r_sign)))) | ((((((fpu___u4___op_div & fpu___rmode_r3[1'h1+:32'h00000001]) & fpu___u4___exp_in_ff) & fpu___u4___op_dn) & ~fpu___u4___r_sign) & (8'h18 > fpu___u4___fi_ldz_2)) & (8'hfe != fpu___u4___exp_out_rnd));
	assign fpu___u4___fract_out_final = ((fpu___u4___inf_out | fpu___u4___ovf0) | fpu_____Vcellinp__u4__output_zero ? 23'h000000 : (fpu___u4___max_num | (fpu___u4___f2i_max & fpu___u4___op_f2i) ? 23'h7fffff : fpu___u4___fract_out_rnd));
	assign fpu___u4___exp_out_final = (((fpu___u4___op_div & fpu___exp_ovf_r[1'h1+:32'h00000001]) & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) | fpu_____Vcellinp__u4__output_zero ? 8'h00 : (((((fpu___u4___op_div & fpu___exp_ovf_r[1'h1+:32'h00000001]) & fpu___exp_ovf_r[1'h0+:32'h00000001]) & fpu___u4___rmode_00) | fpu___u4___inf_out) | (fpu___u4___f2i_max & fpu___u4___op_f2i) ? 8'hff : (fpu___u4___max_num ? 8'hfe : fpu___u4___exp_out_rnd)));
	assign fpu___out_d = {fpu___u4___exp_out_final, fpu___u4___fract_out_final};
	assign fpu___u4___z = (fpu___u4___shft_co | (fpu___exp_ovf_r[1'h1+:32'h00000001] | fpu___u4___exp_in_00)) | ((~fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___u4___exp_in_00) & (fpu___u4___exp_out1_co | fpu___u4___exp_out_00));
	assign fpu___u4___underflow_fmul = ((|fpu___u4___fract_trunc & fpu___u4___z) & ~fpu___u4___exp_in_ff) | ((fpu___u4___fract_out_00 & ~fpu___u4___fract_in_00) & fpu___exp_ovf_r[1'h1+:32'h00000001]);
	assign fpu___u4___undeflow_div = (((~((fpu___exp_ovf_r[1'h1+:32'h00000001] & fpu___exp_ovf_r[1'h0+:32'h00000001]) & fpu___u4___rmode_00) & ~fpu___u4___inf_out) & ~fpu___u4___max_num) & (8'hff != fpu___u4___exp_out_final)) & ((((|fpu___u4___fract_trunc & ~fpu___opb_dn) & ((((((fpu___u4___op_dn & ~fpu___exp_ovf_r[1'h1+:32'h00000001]) & fpu___exp_ovf_r[1'h0+:32'h00000001]) | (fpu___u4___op_dn & fpu___exp_ovf_r[1'h1+:32'h00000001])) | (fpu___u4___op_dn & fpu___u4___div_shft1_co)) | fpu___u4___exp_out_00) | fpu___exp_ovf_r[1'h1+:32'h00000001])) | ((fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) & ((((((fpu___u4___op_dn & (8'h16 < fpu___exp_r)) & (6'h17 > fpu___u4___fi_ldz)) | (((fpu___u4___op_dn & (8'h17 > fpu___exp_r)) & (6'h17 > fpu___u4___fi_ldz)) & ~fpu___remainder_00)) | ((~fpu___u4___op_dn & (fpu___exp_r[3'h7+:32'h00000001] == fpu___u4___exp_div[3'h7+:32'h00000001])) & ~fpu___remainder_00)) | ((~fpu___u4___op_dn & fpu___u4___exp_in_00) & (7'h7f == fpu___u4___exp_div[3'h1+:32'h00000007]))) | ((~fpu___u4___op_dn & (8'h7f > fpu___exp_r)) & (8'h20 < fpu___exp_r))))) | ((~fpu___exp_ovf_r[1'h1+:32'h00000001] & ~fpu___exp_ovf_r[1'h0+:32'h00000001]) & ((((fpu___u4___op_dn & (6'h17 > fpu___u4___fi_ldz)) & fpu___u4___exp_out_00) | (fpu___u4___exp_in_00 & ~fpu___remainder_00)) | ((((~fpu___u4___op_dn & (7'h17 > fpu___u4___ldz_all)) & (8'h01 == fpu___exp_r)) & fpu___u4___exp_out_00) & ~fpu___remainder_00))));
	assign fpu___underflow_d = (fpu___u4___op_div ? fpu___u4___undeflow_div : (fpu___u4___op_mul ? fpu___u4___underflow_fmul : (~fpu___fract_denorm[6'h2f+:32'h00000001] & fpu___u4___exp_out1_co) & ~fpu___u4___dn));
	assign fpu___u4___overflow_fdiv = ((fpu___u4___inf_out | (~fpu___u4___rmode_00 & fpu___u4___max_num)) | ((fpu___exp_r[3'h7+:32'h00000001] & fpu___u4___op_dn) & fpu___u4___exp_out_ff)) | (fpu___exp_ovf_r[1'h0+:32'h00000001] & (fpu___exp_ovf_r[1'h1+:32'h00000001] | fpu___u4___exp_out_ff));
	assign fpu___overflow_d = (fpu___u4___op_div ? fpu___u4___overflow_fdiv : fpu___u4___ovf0 | fpu___u4___ovf1);
	assign fpu___u4___f2i_ine = ((((fpu___u4___f2i_zero & ~fpu___u4___fract_in_00) & ~fpu___opas_r2) | (|fpu___u4___fract_trunc)) | (((fpu___u4___f2i_zero & (8'h80 > fpu___exp_r)) & fpu___opas_r2) & ~fpu___u4___fract_in_00)) | ((fpu___u4___f2i_max & fpu___u4___rmode_11) & (8'h80 > fpu___exp_r));
	assign fpu___ine_d = (fpu___u4___op_f2i ? fpu___u4___f2i_ine : (fpu___u4___op_i2f ? |fpu___u4___fract_trunc : (((fpu___u4___r & ~fpu___u4___dn) | (fpu___u4___s & ~fpu___u4___dn)) | fpu___u4___max_num) | (fpu___u4___op_div & ~fpu___remainder_00)));
endmodule
